module c1355 ( G50gat,G36gat,G29gat,G22gat,G15gat,G8gat,G1gat,G233gat,G227gat,G43gat,G99gat,G71gat,G106gat,G228gat,
G78gat,G226gat,G190gat,G183gat,G169gat,G176gat,G218gat,G211gat,G197gat,G204gat,G64gat,G92gat,G134gat,G232gat,
G162gat,G127gat,G231gat,G155gat,G113gat,G141gat,G229gat,G120gat,G230gat,G85gat,G57gat,G148gat,G225gat,KEYINPUT0,
KEYINPUT1,KEYINPUT2,KEYINPUT3,KEYINPUT4,KEYINPUT5,KEYINPUT6,KEYINPUT7,KEYINPUT8,KEYINPUT9,KEYINPUT10,KEYINPUT11,KEYINPUT12,KEYINPUT13,KEYINPUT14,
KEYINPUT15,KEYINPUT16,KEYINPUT17,KEYINPUT18,KEYINPUT19,KEYINPUT20,KEYINPUT21,KEYINPUT22,KEYINPUT23,KEYINPUT24,KEYINPUT25,KEYINPUT26,KEYINPUT27,KEYINPUT28,
KEYINPUT29,KEYINPUT30,KEYINPUT31,KEYINPUT32,KEYINPUT33,KEYINPUT34,KEYINPUT35,KEYINPUT36,KEYINPUT37,KEYINPUT38,KEYINPUT39,KEYINPUT40,KEYINPUT41,KEYINPUT42,
KEYINPUT43,KEYINPUT44,KEYINPUT45,G1355gat,G1354gat,G1353gat,G1352gat,G1351gat,G1350gat,G1349gat,G1348gat,G1347gat,G1346gat,G1345gat,
G1344gat,G1343gat,G1342gat,G1341gat,G1340gat,G1339gat,G1338gat,G1337gat,G1336gat,G1335gat,G1334gat,G1333gat,G1332gat,G1331gat,
G1330gat,G1329gat,G1328gat,G1327gat,G1326gat,G1325gat,G1324gat );
input G50gat, G36gat, G29gat, G22gat, G15gat, G8gat, G1gat, G233gat,
 G227gat, G43gat, G99gat, G71gat, G106gat, G228gat, G78gat, G226gat, G190gat, G183gat, G169gat, G176gat, G218gat, G211gat,
 G197gat, G204gat, G64gat, G92gat, G134gat, G232gat, G162gat, G127gat, G231gat, G155gat, G113gat, G141gat, G229gat, G120gat,
 G230gat, G85gat, G57gat, G148gat, G225gat, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
 KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
 KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
 KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45;
output G1355gat, G1354gat, G1353gat, G1352gat, G1351gat, G1350gat, G1349gat, G1348gat, G1347gat, G1346gat, G1345gat, G1344gat, G1343gat, G1342gat,
 G1341gat, G1340gat, G1339gat, G1338gat, G1337gat, G1336gat, G1335gat, G1334gat, G1333gat, G1332gat, G1331gat, G1330gat, G1329gat, G1328gat,
 G1327gat, G1326gat, G1325gat, G1324gat;
XOR_X1 U319 ( .A1(w1000), .A2(n287), .ZN(G1355gat) );
NOR_X1 U320 ( .A1(n288), .A2(n289), .ZN(w1001) );
XOR_X1 U321 ( .A1(w1002), .A2(n290), .ZN(G1354gat) );
NOR_X1 U322 ( .A1(n291), .A2(n289), .ZN(w1003) );
XOR_X1 U323 ( .A1(w1004), .A2(n292), .ZN(G1353gat) );
NOR_X1 U324 ( .A1(n293), .A2(n289), .ZN(w1005) );
XOR_X1 U325 ( .A1(w1006), .A2(n294), .ZN(G1352gat) );
NOR_X1 U326 ( .A1(n295), .A2(n289), .ZN(w1007) );
NAND_X1 U327 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(n289) );
XOR_X1 U328 ( .A1(w1008), .A2(n300), .ZN(G1351gat) );
NOR_X1 U329 ( .A1(n288), .A2(n301), .ZN(w1009) );
XOR_X1 U330 ( .A1(w1010), .A2(n302), .ZN(G1350gat) );
NOR_X1 U331 ( .A1(n291), .A2(n301), .ZN(w1011) );
XOR_X1 U332 ( .A1(w1012), .A2(n303), .ZN(G1349gat) );
NOR_X1 U333 ( .A1(n293), .A2(n301), .ZN(w1013) );
XOR_X1 U334 ( .A1(w1014), .A2(n304), .ZN(G1348gat) );
NOR_X1 U335 ( .A1(n295), .A2(n301), .ZN(w1015) );
NAND_X1 U336 ( .A1(n305), .A2(n299), .A3(n306), .A4(n307), .ZN(n301) );
NOR_X1 U337 ( .A1(n308), .A2(n309), .ZN(n307) );
XOR_X1 U338 ( .A1(w1016), .A2(n310), .ZN(G1347gat) );
NOR_X1 U339 ( .A1(n288), .A2(n311), .ZN(w1017) );
XNOR_X1 U340 ( .A1(n312), .A2(n313), .ZN(G1346gat) );
NOR_X1 U341 ( .A1(n291), .A2(n311), .ZN(w1018) );
XOR_X1 U342 ( .A1(w1020), .A2(n314), .ZN(G1345gat) );
NOR_X1 U343 ( .A1(n293), .A2(n311), .ZN(w1021) );
XOR_X1 U344 ( .A1(w1022), .A2(n315), .ZN(G1344gat) );
NOR_X1 U345 ( .A1(n295), .A2(n311), .ZN(w1023) );
NAND_X1 U346 ( .A1(n308), .A2(n299), .A3(n309), .A4(n316), .ZN(n311) );
NOR_X1 U347 ( .A1(n306), .A2(n305), .ZN(n316) );
XOR_X1 U348 ( .A1(w1024), .A2(n317), .ZN(G1343gat) );
NOR_X1 U349 ( .A1(n288), .A2(n318), .ZN(w1025) );
XNOR_X1 U350 ( .A1(n319), .A2(n320), .ZN(G1342gat) );
NOR_X1 U351 ( .A1(n291), .A2(n318), .ZN(w1026) );
XOR_X1 U352 ( .A1(w1028), .A2(n321), .ZN(G1341gat) );
NOR_X1 U353 ( .A1(n293), .A2(n318), .ZN(w1029) );
XOR_X1 U354 ( .A1(w1030), .A2(n322), .ZN(G1340gat) );
NOR_X1 U355 ( .A1(n295), .A2(n318), .ZN(w1031) );
NAND_X1 U356 ( .A1(n323), .A2(n324), .A3(n325), .A4(n299), .ZN(n318) );
NAND_X1 U357 ( .A1(n326), .A2(n327), .ZN(n299) );
OR_X1 U358 ( .A1(n328), .A2(n329), .A3(n330), .ZN(n327) );
OR_X1 U359 ( .A1(n331), .A2(n332), .A3(n333), .ZN(n326) );
XOR_X1 U360 ( .A1(w1032), .A2(n334), .ZN(G1339gat) );
NOR_X1 U361 ( .A1(n325), .A2(n335), .ZN(w1033) );
XOR_X1 U362 ( .A1(w1034), .A2(n336), .ZN(G1338gat) );
NOR_X1 U363 ( .A1(n296), .A2(n335), .ZN(w1035) );
XOR_X1 U364 ( .A1(w1036), .A2(n337), .ZN(G1337gat) );
NOR_X1 U365 ( .A1(n323), .A2(n335), .ZN(w1037) );
XOR_X1 U366 ( .A1(w1038), .A2(n338), .ZN(G1336gat) );
NOR_X1 U367 ( .A1(n298), .A2(n335), .ZN(w1039) );
NAND_X1 U368 ( .A1(n291), .A2(n332), .A3(n295), .A4(n339), .ZN(n335) );
NOR_X1 U369 ( .A1(n288), .A2(n293), .ZN(n332) );
XOR_X1 U370 ( .A1(w1040), .A2(n340), .ZN(G1335gat) );
NOR_X1 U371 ( .A1(n325), .A2(n341), .ZN(w1041) );
XOR_X1 U372 ( .A1(w1042), .A2(n342), .ZN(G1334gat) );
NOR_X1 U373 ( .A1(n296), .A2(n341), .ZN(w1043) );
XOR_X1 U374 ( .A1(w1044), .A2(n343), .ZN(G1333gat) );
NOR_X1 U375 ( .A1(n323), .A2(n341), .ZN(w1045) );
XNOR_X1 U376 ( .A1(n344), .A2(n345), .ZN(G1332gat) );
NOR_X1 U377 ( .A1(n298), .A2(n341), .ZN(n345) );
NAND_X1 U378 ( .A1(n333), .A2(n339), .A3(n330), .A4(n346), .ZN(n341) );
NOR_X1 U379 ( .A1(n328), .A2(n331), .ZN(n346) );
XOR_X1 U380 ( .A1(G50gat), .A2(n347), .ZN(G1331gat) );
NOR_X1 U381 ( .A1(n325), .A2(n348), .ZN(n347) );
XNOR_X1 U382 ( .A1(n349), .A2(n350), .ZN(G1330gat) );
NOR_X1 U383 ( .A1(n296), .A2(n348), .ZN(n350) );
XOR_X1 U384 ( .A1(G36gat), .A2(n351), .ZN(G1329gat) );
NOR_X1 U385 ( .A1(n323), .A2(n348), .ZN(n351) );
XOR_X1 U386 ( .A1(G29gat), .A2(n352), .ZN(G1328gat) );
NOR_X1 U387 ( .A1(n298), .A2(n348), .ZN(n352) );
NAND_X1 U388 ( .A1(n331), .A2(n339), .A3(n328), .A4(n353), .ZN(n348) );
NOR_X1 U389 ( .A1(n333), .A2(n330), .ZN(n353) );
XOR_X1 U390 ( .A1(G22gat), .A2(n354), .ZN(G1327gat) );
NOR_X1 U391 ( .A1(n325), .A2(n355), .ZN(n354) );
XOR_X1 U392 ( .A1(G15gat), .A2(n356), .ZN(G1326gat) );
NOR_X1 U393 ( .A1(n296), .A2(n355), .ZN(n356) );
XOR_X1 U394 ( .A1(G8gat), .A2(n357), .ZN(G1325gat) );
NOR_X1 U395 ( .A1(n323), .A2(n355), .ZN(n357) );
XOR_X1 U396 ( .A1(G1gat), .A2(n358), .ZN(G1324gat) );
NOR_X1 U397 ( .A1(n298), .A2(n355), .ZN(n358) );
NAND_X1 U398 ( .A1(n293), .A2(n329), .A3(n288), .A4(n339), .ZN(n355) );
NAND_X1 U399 ( .A1(n359), .A2(n360), .ZN(n339) );
OR_X1 U400 ( .A1(n308), .A2(n324), .A3(n305), .ZN(n360) );
NOR_X1 U401 ( .A1(n298), .A2(n296), .ZN(n324) );
INV_X1 U402 ( .A1(n306), .ZN(n296) );
OR_X1 U403 ( .A1(n309), .A2(n297), .A3(n306), .ZN(n359) );
XNOR_X1 U404 ( .A1(n361), .A2(n362), .ZN(n306) );
XNOR_X1 U405 ( .A1(G15gat), .A2(n363), .ZN(n362) );
NAND_X1 U406 ( .A1(n364), .A2(n365), .ZN(n363) );
NAND_X1 U407 ( .A1(G233gat), .A2(n366), .A3(G227gat), .ZN(n365) );
XNOR_X1 U408 ( .A1(n367), .A2(n368), .ZN(n366) );
NAND_X1 U409 ( .A1(n369), .A2(n370), .ZN(n364) );
NAND_X1 U410 ( .A1(G227gat), .A2(G233gat), .ZN(n370) );
XNOR_X1 U411 ( .A1(n368), .A2(n371), .ZN(n369) );
XNOR_X1 U412 ( .A1(G43gat), .A2(n372), .ZN(n361) );
XOR_X1 U413 ( .A1(G99gat), .A2(G71gat), .ZN(n372) );
NOR_X1 U414 ( .A1(n323), .A2(n325), .ZN(n297) );
INV_X1 U415 ( .A1(n308), .ZN(n325) );
XNOR_X1 U416 ( .A1(n373), .A2(n374), .ZN(n308) );
XNOR_X1 U417 ( .A1(G106gat), .A2(n375), .ZN(n374) );
NAND_X1 U418 ( .A1(n376), .A2(n377), .ZN(n375) );
NAND_X1 U419 ( .A1(G233gat), .A2(n378), .A3(G228gat), .ZN(n377) );
XNOR_X1 U420 ( .A1(n379), .A2(n380), .ZN(n378) );
NAND_X1 U421 ( .A1(n381), .A2(n382), .ZN(n376) );
NAND_X1 U422 ( .A1(G228gat), .A2(G233gat), .ZN(n382) );
XNOR_X1 U423 ( .A1(n383), .A2(n379), .ZN(n381) );
XNOR_X1 U424 ( .A1(G22gat), .A2(n384), .ZN(n373) );
XOR_X1 U425 ( .A1(G78gat), .A2(G50gat), .ZN(n384) );
INV_X1 U426 ( .A1(n305), .ZN(n323) );
XNOR_X1 U427 ( .A1(n385), .A2(n386), .ZN(n305) );
XNOR_X1 U428 ( .A1(G36gat), .A2(n387), .ZN(n386) );
NAND_X1 U429 ( .A1(n388), .A2(n389), .ZN(n387) );
NAND_X1 U430 ( .A1(G233gat), .A2(n390), .A3(G226gat), .ZN(n389) );
XNOR_X1 U431 ( .A1(n368), .A2(n380), .ZN(n390) );
INV_X1 U432 ( .A1(n383), .ZN(n380) );
NAND_X1 U433 ( .A1(n391), .A2(n392), .ZN(n388) );
NAND_X1 U434 ( .A1(G226gat), .A2(G233gat), .ZN(n392) );
XNOR_X1 U435 ( .A1(n383), .A2(n368), .ZN(n391) );
XNOR_X1 U436 ( .A1(n393), .A2(n394), .ZN(n368) );
XOR_X1 U437 ( .A1(G190gat), .A2(G183gat), .ZN(n394) );
XNOR_X1 U438 ( .A1(G169gat), .A2(G176gat), .ZN(n393) );
XNOR_X1 U439 ( .A1(n395), .A2(n396), .ZN(n383) );
XOR_X1 U440 ( .A1(G218gat), .A2(G211gat), .ZN(n396) );
XNOR_X1 U441 ( .A1(G197gat), .A2(G204gat), .ZN(n395) );
XNOR_X1 U442 ( .A1(G64gat), .A2(n397), .ZN(n385) );
XOR_X1 U443 ( .A1(G92gat), .A2(G8gat), .ZN(n397) );
INV_X1 U444 ( .A1(n328), .ZN(n288) );
XNOR_X1 U445 ( .A1(n398), .A2(n399), .ZN(n328) );
XNOR_X1 U446 ( .A1(G134gat), .A2(n400), .ZN(n399) );
NAND_X1 U447 ( .A1(n401), .A2(n402), .ZN(n400) );
NAND_X1 U448 ( .A1(G233gat), .A2(n403), .A3(G232gat), .ZN(n402) );
XOR_X1 U449 ( .A1(n404), .A2(n405), .ZN(n403) );
NAND_X1 U450 ( .A1(n406), .A2(n407), .ZN(n401) );
NAND_X1 U451 ( .A1(G232gat), .A2(G233gat), .ZN(n407) );
XNOR_X1 U452 ( .A1(n405), .A2(n404), .ZN(n406) );
XNOR_X1 U453 ( .A1(G162gat), .A2(n408), .ZN(n398) );
XOR_X1 U454 ( .A1(G218gat), .A2(G190gat), .ZN(n408) );
NOR_X1 U455 ( .A1(n295), .A2(n291), .ZN(n329) );
INV_X1 U456 ( .A1(n333), .ZN(n291) );
XNOR_X1 U457 ( .A1(n409), .A2(n410), .ZN(n333) );
XNOR_X1 U458 ( .A1(G127gat), .A2(n411), .ZN(n410) );
NAND_X1 U459 ( .A1(n412), .A2(n413), .ZN(n411) );
NAND_X1 U460 ( .A1(G231gat), .A2(n414), .A3(G233gat), .ZN(n413) );
XNOR_X1 U461 ( .A1(n415), .A2(n416), .ZN(n414) );
NAND_X1 U462 ( .A1(n417), .A2(n418), .ZN(n412) );
NAND_X1 U463 ( .A1(G233gat), .A2(G231gat), .ZN(n418) );
XNOR_X1 U464 ( .A1(n419), .A2(n415), .ZN(n417) );
XNOR_X1 U465 ( .A1(G155gat), .A2(n420), .ZN(n409) );
XOR_X1 U466 ( .A1(G211gat), .A2(G183gat), .ZN(n420) );
INV_X1 U467 ( .A1(n331), .ZN(n295) );
NAND_X1 U468 ( .A1(n421), .A2(n422), .ZN(n331) );
NAND_X1 U469 ( .A1(n423), .A2(n424), .ZN(n422) );
NAND_X1 U470 ( .A1(n425), .A2(n426), .ZN(n424) );
NAND_X1 U471 ( .A1(n425), .A2(n426), .A3(n427), .ZN(n421) );
INV_X1 U472 ( .A1(n423), .ZN(n427) );
XNOR_X1 U473 ( .A1(n428), .A2(n429), .ZN(n423) );
XOR_X1 U474 ( .A1(G197gat), .A2(G169gat), .ZN(n429) );
XNOR_X1 U475 ( .A1(G113gat), .A2(G141gat), .ZN(n428) );
NAND_X1 U476 ( .A1(n430), .A2(n431), .ZN(n426) );
NAND_X1 U477 ( .A1(G229gat), .A2(G233gat), .ZN(n431) );
XNOR_X1 U478 ( .A1(n419), .A2(n405), .ZN(n430) );
NAND_X1 U479 ( .A1(G233gat), .A2(n432), .A3(G229gat), .ZN(n425) );
XNOR_X1 U480 ( .A1(n405), .A2(n416), .ZN(n432) );
INV_X1 U481 ( .A1(n419), .ZN(n416) );
XNOR_X1 U482 ( .A1(n433), .A2(n434), .ZN(n419) );
XOR_X1 U483 ( .A1(G8gat), .A2(G22gat), .ZN(n434) );
XNOR_X1 U484 ( .A1(G15gat), .A2(G1gat), .ZN(n433) );
XNOR_X1 U485 ( .A1(n435), .A2(n436), .ZN(n405) );
XNOR_X1 U486 ( .A1(G50gat), .A2(n349), .ZN(n436) );
INV_X1 U487 ( .A1(G43gat), .ZN(n349) );
XNOR_X1 U488 ( .A1(G29gat), .A2(G36gat), .ZN(n435) );
INV_X1 U489 ( .A1(n330), .ZN(n293) );
XNOR_X1 U490 ( .A1(n437), .A2(n438), .ZN(n330) );
XNOR_X1 U491 ( .A1(G120gat), .A2(n439), .ZN(n438) );
NAND_X1 U492 ( .A1(n440), .A2(n441), .ZN(n439) );
NAND_X1 U493 ( .A1(G233gat), .A2(n442), .A3(G230gat), .ZN(n441) );
XOR_X1 U494 ( .A1(n404), .A2(n415), .ZN(n442) );
NAND_X1 U495 ( .A1(n443), .A2(n444), .ZN(n440) );
NAND_X1 U496 ( .A1(G230gat), .A2(G233gat), .ZN(n444) );
XNOR_X1 U497 ( .A1(n415), .A2(n404), .ZN(n443) );
XNOR_X1 U498 ( .A1(n445), .A2(n446), .ZN(n404) );
XOR_X1 U499 ( .A1(G99gat), .A2(G92gat), .ZN(n446) );
XNOR_X1 U500 ( .A1(G106gat), .A2(G85gat), .ZN(n445) );
XNOR_X1 U501 ( .A1(n447), .A2(n448), .ZN(n415) );
XOR_X1 U502 ( .A1(G78gat), .A2(G71gat), .ZN(n448) );
XNOR_X1 U503 ( .A1(G57gat), .A2(G64gat), .ZN(n447) );
XNOR_X1 U504 ( .A1(G148gat), .A2(n449), .ZN(n437) );
XOR_X1 U505 ( .A1(G204gat), .A2(G176gat), .ZN(n449) );
INV_X1 U506 ( .A1(n309), .ZN(n298) );
NAND_X1 U507 ( .A1(n450), .A2(n451), .ZN(n309) );
NAND_X1 U508 ( .A1(n452), .A2(n453), .ZN(n451) );
NAND_X1 U509 ( .A1(n454), .A2(n455), .ZN(n453) );
NAND_X1 U510 ( .A1(n454), .A2(n455), .A3(n456), .ZN(n450) );
INV_X1 U511 ( .A1(n452), .ZN(n456) );
XNOR_X1 U512 ( .A1(n457), .A2(n458), .ZN(n452) );
XNOR_X1 U513 ( .A1(G85gat), .A2(n344), .ZN(n458) );
INV_X1 U514 ( .A1(G57gat), .ZN(n344) );
XNOR_X1 U515 ( .A1(G1gat), .A2(G29gat), .ZN(n457) );
NAND_X1 U516 ( .A1(n459), .A2(n460), .ZN(n455) );
NAND_X1 U517 ( .A1(G225gat), .A2(G233gat), .ZN(n460) );
XNOR_X1 U518 ( .A1(n371), .A2(n379), .ZN(n459) );
NAND_X1 U519 ( .A1(G233gat), .A2(n461), .A3(G225gat), .ZN(n454) );
XNOR_X1 U520 ( .A1(n379), .A2(n367), .ZN(n461) );
INV_X1 U521 ( .A1(n371), .ZN(n367) );
XNOR_X1 U522 ( .A1(n462), .A2(n463), .ZN(n371) );
XNOR_X1 U523 ( .A1(G134gat), .A2(n319), .ZN(n463) );
INV_X1 U524 ( .A1(G127gat), .ZN(w1027) );
XNOR_X1 U525 ( .A1(G113gat), .A2(G120gat), .ZN(n462) );
XNOR_X1 U526 ( .A1(n464), .A2(n465), .ZN(n379) );
XNOR_X1 U527 ( .A1(G162gat), .A2(n312), .ZN(n465) );
INV_X1 U528 ( .A1(G155gat), .ZN(w1019) );
XNOR_X1 U529 ( .A1(G141gat), .A2(G148gat), .ZN(n464) );
XOR_X1 X1000 ( .A1(G218gat), .A2(KEYINPUT0), .ZN(w1000) );
XNOR_X1 X1001 ( .A1(w1001), .A2(KEYINPUT1), .ZN(n287) );
XOR_X1 X1002 ( .A1(G211gat), .A2(KEYINPUT2), .ZN(w1002) );
XNOR_X1 X1003 ( .A1(w1003), .A2(KEYINPUT3), .ZN(n290) );
XOR_X1 X1004 ( .A1(G204gat), .A2(KEYINPUT4), .ZN(w1004) );
XNOR_X1 X1005 ( .A1(w1005), .A2(KEYINPUT5), .ZN(n292) );
XOR_X1 X1006 ( .A1(G197gat), .A2(KEYINPUT6), .ZN(w1006) );
XNOR_X1 X1007 ( .A1(w1007), .A2(KEYINPUT7), .ZN(n294) );
XOR_X1 X1008 ( .A1(G190gat), .A2(KEYINPUT8), .ZN(w1008) );
XNOR_X1 X1009 ( .A1(w1009), .A2(KEYINPUT9), .ZN(n300) );
XOR_X1 X1010 ( .A1(G183gat), .A2(KEYINPUT10), .ZN(w1010) );
XNOR_X1 X1011 ( .A1(w1011), .A2(KEYINPUT11), .ZN(n302) );
XOR_X1 X1012 ( .A1(G176gat), .A2(KEYINPUT12), .ZN(w1012) );
XNOR_X1 X1013 ( .A1(w1013), .A2(KEYINPUT13), .ZN(n303) );
XOR_X1 X1014 ( .A1(G169gat), .A2(KEYINPUT14), .ZN(w1014) );
XNOR_X1 X1015 ( .A1(w1015), .A2(KEYINPUT15), .ZN(n304) );
XOR_X1 X1016 ( .A1(G162gat), .A2(KEYINPUT16), .ZN(w1016) );
XNOR_X1 X1017 ( .A1(w1017), .A2(KEYINPUT17), .ZN(n310) );
XOR_X1 X1018 ( .A1(w1018), .A2(KEYINPUT18), .ZN(n313) );
XNOR_X1 X1019 ( .A1(w1019), .A2(KEYINPUT19), .ZN(n312) );
XOR_X1 X1020 ( .A1(G148gat), .A2(KEYINPUT20), .ZN(w1020) );
XNOR_X1 X1021 ( .A1(w1021), .A2(KEYINPUT21), .ZN(n314) );
XOR_X1 X1022 ( .A1(G141gat), .A2(KEYINPUT22), .ZN(w1022) );
XNOR_X1 X1023 ( .A1(w1023), .A2(KEYINPUT23), .ZN(n315) );
XOR_X1 X1024 ( .A1(G134gat), .A2(KEYINPUT24), .ZN(w1024) );
XNOR_X1 X1025 ( .A1(w1025), .A2(KEYINPUT25), .ZN(n317) );
XOR_X1 X1026 ( .A1(w1026), .A2(KEYINPUT26), .ZN(n320) );
XNOR_X1 X1027 ( .A1(w1027), .A2(KEYINPUT27), .ZN(n319) );
XOR_X1 X1028 ( .A1(G120gat), .A2(KEYINPUT28), .ZN(w1028) );
XNOR_X1 X1029 ( .A1(w1029), .A2(KEYINPUT29), .ZN(n321) );
XOR_X1 X1030 ( .A1(G113gat), .A2(KEYINPUT30), .ZN(w1030) );
XNOR_X1 X1031 ( .A1(w1031), .A2(KEYINPUT31), .ZN(n322) );
XOR_X1 X1032 ( .A1(G106gat), .A2(KEYINPUT32), .ZN(w1032) );
XNOR_X1 X1033 ( .A1(w1033), .A2(KEYINPUT33), .ZN(n334) );
XOR_X1 X1034 ( .A1(G99gat), .A2(KEYINPUT34), .ZN(w1034) );
XNOR_X1 X1035 ( .A1(w1035), .A2(KEYINPUT35), .ZN(n336) );
XOR_X1 X1036 ( .A1(G92gat), .A2(KEYINPUT36), .ZN(w1036) );
XNOR_X1 X1037 ( .A1(w1037), .A2(KEYINPUT37), .ZN(n337) );
XOR_X1 X1038 ( .A1(G85gat), .A2(KEYINPUT38), .ZN(w1038) );
XNOR_X1 X1039 ( .A1(w1039), .A2(KEYINPUT39), .ZN(n338) );
XOR_X1 X1040 ( .A1(G78gat), .A2(KEYINPUT40), .ZN(w1040) );
XNOR_X1 X1041 ( .A1(w1041), .A2(KEYINPUT41), .ZN(n340) );
XOR_X1 X1042 ( .A1(G71gat), .A2(KEYINPUT42), .ZN(w1042) );
XNOR_X1 X1043 ( .A1(w1043), .A2(KEYINPUT43), .ZN(n342) );
XOR_X1 X1044 ( .A1(G64gat), .A2(KEYINPUT44), .ZN(w1044) );
XNOR_X1 X1045 ( .A1(w1045), .A2(KEYINPUT45), .ZN(n343) );
