module c2670 ( G2066,G1083,G452,G1986,G1981,G1976,G8,G1956,G2072,G1341,G2067,G1996,G40,G1384,
G868,G2,G15,G661,G108,G57,G120,G69,G567,G1971,G142,G106,G130,G118,
G14,G37,G96,G82,G132,G44,G2106,G7,G3,G1,G36,G483,G94,G2090,
G2084,G2078,G2100,G11,G29,G28,G138,G102,G126,G114,G1991,G141,G105,G129,
G117,G135,G99,G123,G111,G131,G95,G119,G107,G137,G101,G125,G113,G136,
G100,G124,G112,G139,G103,G127,G115,G140,G2104,G2105,G104,G128,G116,G16,
G89,G76,G51,G63,G1348,G49,G87,G74,G651,G85,G72,G47,G60,G90,
G77,G52,G64,G91,G78,G53,G65,G88,G75,G50,G62,G86,G73,G48,
G61,G23,G22,G19,G20,G4,G5,G1961,G21,G1966,G93,G80,G55,G67,
G559,G860,G92,G79,G54,G66,G81,G543,G68,G43,G56,KEYINPUT0,KEYINPUT1,KEYINPUT2,
KEYINPUT3,KEYINPUT4,KEYINPUT5,KEYINPUT6,KEYINPUT7,KEYINPUT8,KEYINPUT9,KEYINPUT10,KEYINPUT11,KEYINPUT12,KEYINPUT13,G2678,KEYINPUT14,KEYINPUT15,
G2096,KEYINPUT16,KEYINPUT17,KEYINPUT18,KEYINPUT19,KEYINPUT20,KEYINPUT21,KEYINPUT22,KEYINPUT23,KEYINPUT24,KEYINPUT25,KEYINPUT26,KEYINPUT27,G2474,
KEYINPUT28,KEYINPUT29,KEYINPUT30,KEYINPUT31,KEYINPUT32,KEYINPUT33,KEYINPUT34,KEYINPUT35,KEYINPUT36,KEYINPUT37,KEYINPUT38,KEYINPUT39,KEYINPUT40,KEYINPUT41,
KEYINPUT42,KEYINPUT43,KEYINPUT44,KEYINPUT45,KEYINPUT46,KEYINPUT47,KEYINPUT48,KEYINPUT49,KEYINPUT50,KEYINPUT51,KEYINPUT52,KEYINPUT53,G2430,KEYINPUT54,
G2427,KEYINPUT55,KEYINPUT56,KEYINPUT57,KEYINPUT58,KEYINPUT59,KEYINPUT60,KEYINPUT61,G2446,KEYINPUT62,G2443,KEYINPUT63,G2454,KEYINPUT64,
G2451,KEYINPUT65,KEYINPUT66,KEYINPUT67,G2438,KEYINPUT68,G2435,KEYINPUT69,KEYINPUT70,KEYINPUT71,KEYINPUT72,KEYINPUT73,KEYINPUT74,KEYINPUT75,
KEYINPUT76,KEYINPUT77,KEYINPUT78,KEYINPUT79,KEYINPUT80,KEYINPUT81,KEYINPUT82,KEYINPUT83,KEYINPUT84,KEYINPUT85,KEYINPUT86,KEYINPUT87,KEYINPUT88,KEYINPUT89,
G27,KEYINPUT90,KEYINPUT91,G34,KEYINPUT92,KEYINPUT93,G35,KEYINPUT94,KEYINPUT95,G25,KEYINPUT96,KEYINPUT97,G32,KEYINPUT98,
KEYINPUT99,G26,KEYINPUT100,KEYINPUT101,G33,KEYINPUT102,KEYINPUT103,KEYINPUT104,KEYINPUT105,KEYINPUT106,KEYINPUT107,KEYINPUT108,KEYINPUT109,KEYINPUT110,
KEYINPUT111,KEYINPUT112,KEYINPUT113,KEYINPUT114,KEYINPUT115,KEYINPUT116,KEYINPUT117,KEYINPUT118,KEYINPUT119,KEYINPUT120,KEYINPUT121,KEYINPUT122,KEYINPUT123,KEYINPUT124,
KEYINPUT125,KEYINPUT126,KEYINPUT127,KEYINPUT128,G24,KEYINPUT129,KEYINPUT130,G6,KEYINPUT131,G231,G331,G323,G280,G321,
G337,G411,G384,G369,G367,G409,G335,G350,G391,G401,G397,G395,G329,G311,
G308,G297,G295,G284,G282,G261,G325,G259,G238,G237,G236,G235,G234,G225,
G227,G229,G221,G220,G219,G218,G217,G223,G188,G176,G319,G173,G171,G168,
G164,G158,G156,G153,G150,G160,G162,G286,G288,G290,G301,G299,G166,G303,
G305,G148,G145 );
input G2066, G1083, G452, G1986, G1981, G1976, G8, G1956, G2072, G1341, G2067, G1996,
 G40, G1384, G868, G2, G15, G661, G108, G57, G120, G69, G567, G1971, G142, G106,
 G130, G118, G14, G37, G96, G82, G132, G44, G2106, G7, G3, G1, G36, G483,
 G94, G2090, G2084, G2078, G2100, G11, G29, G28, G138, G102, G126, G114, G1991, G141,
 G105, G129, G117, G135, G99, G123, G111, G131, G95, G119, G107, G137, G101, G125,
 G113, G136, G100, G124, G112, G139, G103, G127, G115, G140, G2104, G2105, G104, G128,
 G116, G16, G89, G76, G51, G63, G1348, G49, G87, G74, G651, G85, G72, G47,
 G60, G90, G77, G52, G64, G91, G78, G53, G65, G88, G75, G50, G62, G86,
 G73, G48, G61, G23, G22, G19, G20, G4, G5, G1961, G21, G1966, G93, G80,
 G55, G67, G559, G860, G92, G79, G54, G66, G81, G543, G68, G43, G56, KEYINPUT0,
 KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, G2678,
 KEYINPUT14, KEYINPUT15, G2096, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
 KEYINPUT27, G2474, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39,
 KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
 G2430, KEYINPUT54, G2427, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, G2446, KEYINPUT62, G2443, KEYINPUT63,
 G2454, KEYINPUT64, G2451, KEYINPUT65, KEYINPUT66, KEYINPUT67, G2438, KEYINPUT68, G2435, KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73,
 KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
 KEYINPUT88, KEYINPUT89, G27, KEYINPUT90, KEYINPUT91, G34, KEYINPUT92, KEYINPUT93, G35, KEYINPUT94, KEYINPUT95, G25, KEYINPUT96, KEYINPUT97,
 G32, KEYINPUT98, KEYINPUT99, G26, KEYINPUT100, KEYINPUT101, G33, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
 KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122,
 KEYINPUT123, KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT128, G24, KEYINPUT129, KEYINPUT130, G6, KEYINPUT131;
output G231, G331, G323, G280, G321, G337, G411, G384, G369, G367, G409, G335, G350, G391,
 G401, G397, G395, G329, G311, G308, G297, G295, G284, G282, G261, G325, G259, G238,
 G237, G236, G235, G234, G225, G227, G229, G221, G220, G219, G218, G217, G223, G188,
 G176, G319, G173, G171, G168, G164, G158, G156, G153, G150, G160, G162, G286, G288,
 G290, G301, G299, G166, G303, G305, G148, G145;
INV_X1 U437 ( .A1(1'b1), .ZN(G231) );
BUF_X1 U439 ( .A1(G295), .ZN(G331) );
BUF_X1 U440 ( .A1(G282), .ZN(G323) );
BUF_X1 U441 ( .A1(G297), .ZN(G280) );
BUF_X1 U442 ( .A1(G284), .ZN(G321) );
INV_X1 U443 ( .A1(G2066), .ZN(n414) );
INV_X1 U444 ( .A1(n414), .ZN(G337) );
INV_X1 U445 ( .A1(n414), .ZN(G411) );
INV_X1 U446 ( .A1(n414), .ZN(G384) );
BUF_X1 U447 ( .A1(G1083), .ZN(G369) );
BUF_X1 U448 ( .A1(G1083), .ZN(G367) );
INV_X1 U449 ( .A1(G452), .ZN(n420) );
INV_X1 U450 ( .A1(n420), .ZN(G409) );
INV_X1 U451 ( .A1(n420), .ZN(G335) );
INV_X1 U452 ( .A1(n420), .ZN(G350) );
INV_X1 U453 ( .A1(n420), .ZN(G391) );
INV_X1 U454 ( .A1(n425), .ZN(G401) );
INV_X1 U455 ( .A1(n426), .ZN(G397) );
INV_X1 U456 ( .A1(n427), .ZN(G395) );
NAND_X1 U457 ( .A1(n428), .A2(n429), .A3(n430), .ZN(G329) );
OR_X1 U458 ( .A1(n431), .A2(n432), .ZN(n430) );
NAND_X1 U459 ( .A1(n433), .A2(n434), .ZN(n429) );
NAND_X1 U460 ( .A1(n435), .A2(n436), .ZN(n433) );
NAND_X1 U461 ( .A1(n432), .A2(n437), .ZN(n436) );
INV_X1 U462 ( .A1(n438), .ZN(n435) );
NAND_X1 U463 ( .A1(n437), .A2(n438), .ZN(n428) );
NAND_X1 U464 ( .A1(n431), .A2(n439), .ZN(n438) );
NAND_X1 U465 ( .A1(n440), .A2(n441), .A3(n432), .ZN(n439) );
NAND_X1 U466 ( .A1(n442), .A2(n443), .ZN(n431) );
NAND_X1 U467 ( .A1(n444), .A2(n445), .ZN(n443) );
NAND_X1 U468 ( .A1(n446), .A2(n447), .A3(n448), .A4(n449), .ZN(n445) );
NAND_X1 U469 ( .A1(n432), .A2(G290), .A3(G1986), .ZN(n449) );
NAND_X1 U470 ( .A1(G1981), .A2(n450), .ZN(n448) );
NAND_X1 U471 ( .A1(n451), .A2(n452), .ZN(n450) );
NAND_X1 U472 ( .A1(n453), .A2(G305), .ZN(n452) );
NAND_X1 U473 ( .A1(n454), .A2(G305), .ZN(n447) );
INV_X1 U474 ( .A1(n451), .ZN(n454) );
NAND_X1 U475 ( .A1(n455), .A2(n456), .ZN(n451) );
OR_X1 U476 ( .A1(G288), .A2(G1976), .ZN(n455) );
NAND_X1 U477 ( .A1(n456), .A2(n457), .ZN(n446) );
NAND_X1 U478 ( .A1(n458), .A2(n459), .A3(n460), .ZN(n456) );
OR_X1 U479 ( .A1(n461), .A2(n457), .ZN(n460) );
NAND_X1 U480 ( .A1(n462), .A2(n463), .A3(n464), .ZN(n459) );
INV_X1 U481 ( .A1(n465), .ZN(n464) );
NAND_X1 U482 ( .A1(n466), .A2(G303), .A3(G8), .ZN(n458) );
NAND_X1 U483 ( .A1(n465), .A2(n467), .ZN(n466) );
NAND_X1 U484 ( .A1(n462), .A2(n463), .ZN(n467) );
NAND_X1 U485 ( .A1(n468), .A2(n469), .A3(n470), .ZN(n463) );
OR_X1 U486 ( .A1(n471), .A2(G171), .ZN(n470) );
NAND_X1 U487 ( .A1(G8), .A2(G286), .A3(n472), .ZN(n469) );
INV_X1 U488 ( .A1(n473), .ZN(n472) );
NAND_X1 U489 ( .A1(n474), .A2(n475), .A3(n476), .ZN(n468) );
NAND_X1 U490 ( .A1(n471), .A2(G171), .ZN(n476) );
NAND_X1 U491 ( .A1(n477), .A2(n478), .ZN(n471) );
NAND_X1 U492 ( .A1(n479), .A2(n480), .A3(n481), .ZN(n478) );
NAND_X1 U493 ( .A1(G1956), .A2(n482), .ZN(n480) );
NAND_X1 U494 ( .A1(G2072), .A2(n483), .ZN(n479) );
NAND_X1 U495 ( .A1(n484), .A2(n485), .A3(n486), .ZN(n477) );
NAND_X1 U496 ( .A1(n487), .A2(n482), .ZN(n485) );
NAND_X1 U497 ( .A1(n488), .A2(n489), .A3(n490), .ZN(n487) );
NAND_X1 U498 ( .A1(G1956), .A2(G299), .ZN(n490) );
NAND_X1 U499 ( .A1(G1341), .A2(n491), .ZN(n489) );
OR_X1 U500 ( .A1(n492), .A2(n493), .ZN(n488) );
NAND_X1 U501 ( .A1(n483), .A2(n494), .ZN(n484) );
NAND_X1 U502 ( .A1(n495), .A2(n496), .A3(n497), .ZN(n494) );
NAND_X1 U503 ( .A1(G2072), .A2(G299), .ZN(n497) );
NAND_X1 U504 ( .A1(G2067), .A2(n498), .ZN(n496) );
NAND_X1 U505 ( .A1(n493), .A2(n441), .ZN(n498) );
NAND_X1 U506 ( .A1(G1996), .A2(n499), .ZN(n495) );
NAND_X1 U507 ( .A1(n483), .A2(n500), .ZN(n475) );
NAND_X1 U508 ( .A1(n482), .A2(n501), .ZN(n474) );
NAND_X1 U509 ( .A1(n473), .A2(G168), .ZN(n462) );
NAND_X1 U510 ( .A1(n502), .A2(n503), .ZN(n473) );
NAND_X1 U511 ( .A1(G8), .A2(n504), .A3(n483), .ZN(n503) );
NAND_X1 U512 ( .A1(n453), .A2(n505), .ZN(n502) );
NAND_X1 U513 ( .A1(n506), .A2(n507), .ZN(n465) );
NAND_X1 U514 ( .A1(G8), .A2(n508), .A3(n483), .ZN(n507) );
INV_X1 U515 ( .A1(n482), .ZN(n483) );
NAND_X1 U516 ( .A1(n453), .A2(n509), .ZN(n506) );
INV_X1 U517 ( .A1(n457), .ZN(n453) );
NAND_X1 U518 ( .A1(G8), .A2(n482), .ZN(n457) );
NAND_X1 U519 ( .A1(G40), .A2(G160), .A3(n510), .A4(n511), .ZN(n482) );
NAND_X1 U520 ( .A1(n432), .A2(n512), .ZN(n444) );
NAND_X1 U521 ( .A1(n513), .A2(n514), .ZN(n512) );
OR_X1 U522 ( .A1(G290), .A2(G1986), .ZN(n514) );
NAND_X1 U523 ( .A1(n432), .A2(n515), .ZN(n442) );
AND_X1 U524 ( .A1(G160), .A2(n516), .A3(G40), .ZN(n432) );
NAND_X1 U525 ( .A1(n510), .A2(n511), .ZN(n516) );
INV_X1 U526 ( .A1(G1384), .ZN(n511) );
INV_X1 U527 ( .A1(G150), .ZN(G311) );
INV_X1 U528 ( .A1(G225), .ZN(G308) );
NAND_X1 U529 ( .A1(n517), .A2(n518), .ZN(G297) );
NAND_X1 U530 ( .A1(G868), .A2(G286), .ZN(n518) );
NAND_X1 U531 ( .A1(G299), .A2(n519), .ZN(n517) );
NAND_X1 U532 ( .A1(n520), .A2(n521), .ZN(G295) );
NAND_X1 U533 ( .A1(n522), .A2(n519), .ZN(n521) );
NAND_X1 U534 ( .A1(G868), .A2(n523), .ZN(w1000) );
XNOR_X1 U535 ( .A1(n524), .A2(n525), .ZN(w1074) );
XNOR_X1 U536 ( .A1(n526), .A2(n527), .ZN(w1080) );
NAND_X1 U537 ( .A1(n528), .A2(n529), .ZN(G284) );
NAND_X1 U538 ( .A1(G868), .A2(G301), .ZN(n529) );
NAND_X1 U539 ( .A1(n499), .A2(n519), .ZN(n528) );
NAND_X1 U540 ( .A1(n530), .A2(n531), .ZN(G282) );
NAND_X1 U541 ( .A1(G868), .A2(n526), .ZN(n531) );
NAND_X1 U542 ( .A1(n532), .A2(n519), .ZN(n530) );
INV_X1 U543 ( .A1(G868), .ZN(n519) );
INV_X1 U544 ( .A1(G325), .ZN(G261) );
NOR_X1 U545 ( .A1(n533), .A2(n534), .ZN(G325) );
NAND_X1 U546 ( .A1(G2), .A2(G15), .A3(G661), .ZN(G259) );
INV_X1 U547 ( .A1(G108), .ZN(G238) );
INV_X1 U548 ( .A1(G57), .ZN(G237) );
INV_X1 U549 ( .A1(G120), .ZN(G236) );
INV_X1 U550 ( .A1(G69), .ZN(G235) );
NAND_X1 U551 ( .A1(G567), .A2(n535), .ZN(G234) );
NAND_X1 U552 ( .A1(n426), .A2(n425), .A3(n427), .A4(n536), .ZN(G225) );
NOR_X1 U553 ( .A1(n537), .A2(G229), .A3(G227), .ZN(w1018) );
XOR_X1 U554 ( .A1(n538), .A2(n539), .ZN(w1012) );
XOR_X1 U555 ( .A1(n540), .A2(n541), .ZN(w1011) );
XNOR_X1 U556 ( .A1(w1008), .A2(n434), .ZN(w1007) );
XNOR_X1 U557 ( .A1(n504), .A2(w1010), .ZN(n540) );
XOR_X1 U558 ( .A1(n542), .A2(n543), .ZN(w1015) );
XNOR_X1 U559 ( .A1(w1014), .A2(n544), .ZN(w1013) );
XNOR_X1 U560 ( .A1(w1016), .A2(w1017), .ZN(n542) );
XOR_X1 U561 ( .A1(n545), .A2(n546), .ZN(w1022) );
XOR_X1 U562 ( .A1(w1020), .A2(w1021), .ZN(w1019) );
XOR_X1 U563 ( .A1(n547), .A2(n548), .ZN(w1030) );
XOR_X1 U564 ( .A1(n549), .A2(n550), .ZN(w1029) );
XNOR_X1 U565 ( .A1(n551), .A2(w1026), .ZN(w1025) );
XNOR_X1 U566 ( .A1(w1028), .A2(n441), .ZN(n549) );
XOR_X1 U567 ( .A1(n552), .A2(n553), .ZN(w1033) );
XNOR_X1 U568 ( .A1(n509), .A2(w1032), .ZN(w1031) );
INV_X1 U569 ( .A1(G1971), .ZN(n509) );
XNOR_X1 U570 ( .A1(w1034), .A2(w1035), .ZN(n552) );
NAND_X1 U571 ( .A1(n554), .A2(n555), .ZN(w1036) );
XOR_X1 U572 ( .A1(n556), .A2(n557), .ZN(w1038) );
XOR_X1 U573 ( .A1(n558), .A2(n559), .ZN(w1046) );
XOR_X1 U574 ( .A1(n560), .A2(n561), .ZN(w1044) );
XNOR_X1 U575 ( .A1(G162), .A2(n562), .ZN(w1041) );
XNOR_X1 U576 ( .A1(n563), .A2(G164), .ZN(n560) );
XOR_X1 U577 ( .A1(n564), .A2(n565), .ZN(w1050) );
XNOR_X1 U578 ( .A1(n440), .A2(n566), .ZN(w1047) );
XNOR_X1 U579 ( .A1(n567), .A2(n568), .ZN(n564) );
NAND_X1 U580 ( .A1(n569), .A2(n570), .A3(n571), .A4(n572), .ZN(w1051) );
NAND_X1 U581 ( .A1(G142), .A2(n573), .ZN(n572) );
NAND_X1 U582 ( .A1(G106), .A2(n574), .ZN(n571) );
NAND_X1 U583 ( .A1(G130), .A2(n575), .ZN(n570) );
NAND_X1 U584 ( .A1(G118), .A2(n576), .ZN(n569) );
NAND_X1 U585 ( .A1(n577), .A2(G14), .ZN(w1052) );
XOR_X1 U586 ( .A1(n578), .A2(n579), .ZN(w1056) );
XOR_X1 U587 ( .A1(w1054), .A2(w1055), .ZN(w1053) );
XNOR_X1 U588 ( .A1(n580), .A2(n492), .ZN(w1058) );
XOR_X1 U589 ( .A1(n581), .A2(n582), .ZN(w1067) );
XOR_X1 U590 ( .A1(n583), .A2(n584), .ZN(w1059) );
XNOR_X1 U591 ( .A1(w1062), .A2(w1063), .ZN(w1061) );
XNOR_X1 U592 ( .A1(w1064), .A2(w1065), .ZN(n583) );
XOR_X1 U593 ( .A1(n585), .A2(w1066), .ZN(n581) );
XNOR_X1 U594 ( .A1(w1068), .A2(w1069), .ZN(n585) );
NAND_X1 U595 ( .A1(n586), .A2(n555), .ZN(w1070) );
INV_X1 U596 ( .A1(G37), .ZN(n555) );
XOR_X1 U597 ( .A1(n587), .A2(n588), .ZN(w1086) );
XNOR_X1 U598 ( .A1(n527), .A2(n589), .ZN(w1081) );
INV_X1 U599 ( .A1(n524), .ZN(w1075) );
XNOR_X1 U600 ( .A1(n590), .A2(n591), .ZN(w1078) );
XNOR_X1 U601 ( .A1(n481), .A2(n499), .ZN(n591) );
INV_X1 U602 ( .A1(G299), .ZN(w1077) );
XNOR_X1 U603 ( .A1(n532), .A2(n522), .ZN(n590) );
XNOR_X1 U604 ( .A1(n592), .A2(n593), .ZN(w1084) );
XNOR_X1 U605 ( .A1(G166), .A2(G288), .ZN(n593) );
XNOR_X1 U606 ( .A1(G290), .A2(G305), .ZN(n592) );
XNOR_X1 U607 ( .A1(G168), .A2(G171), .ZN(n587) );
INV_X1 U608 ( .A1(G96), .ZN(G221) );
INV_X1 U609 ( .A1(G82), .ZN(G220) );
INV_X1 U610 ( .A1(G132), .ZN(G219) );
INV_X1 U611 ( .A1(G44), .ZN(G218) );
NAND_X1 U612 ( .A1(G2106), .A2(n535), .ZN(G217) );
INV_X1 U613 ( .A1(G223), .ZN(n535) );
NAND_X1 U614 ( .A1(G7), .A2(G661), .ZN(G223) );
NAND_X1 U615 ( .A1(n594), .A2(n595), .ZN(G188) );
NAND_X1 U616 ( .A1(G3), .A2(G1), .ZN(n595) );
NAND_X1 U617 ( .A1(G36), .A2(n594), .ZN(G176) );
AND_X1 U618 ( .A1(G661), .A2(G319), .A3(G483), .ZN(n594) );
INV_X1 U619 ( .A1(n537), .ZN(G319) );
NAND_X1 U620 ( .A1(n596), .A2(n597), .ZN(n537) );
NAND_X1 U621 ( .A1(G2106), .A2(n534), .ZN(n597) );
NAND_X1 U622 ( .A1(G44), .A2(G132), .A3(G82), .A4(G96), .ZN(n534) );
NAND_X1 U623 ( .A1(G567), .A2(n533), .ZN(n596) );
NAND_X1 U624 ( .A1(G69), .A2(G120), .A3(G57), .A4(G108), .ZN(n533) );
AND_X1 U625 ( .A1(G94), .A2(G452), .ZN(G173) );
INV_X1 U626 ( .A1(G301), .ZN(w1087) );
INV_X1 U627 ( .A1(G286), .ZN(G168) );
INV_X1 U628 ( .A1(n510), .ZN(w1045) );
NAND_X1 U629 ( .A1(G2090), .A2(G2084), .A3(G2078), .A4(G2072), .ZN(G158) );
NAND_X1 U630 ( .A1(n598), .A2(n544), .ZN(w1089) );
INV_X1 U631 ( .A1(G2100), .ZN(n544) );
XOR_X1 U632 ( .A1(n556), .A2(w1088), .ZN(n598) );
OR_X1 U633 ( .A1(n599), .A2(n532), .ZN(G153) );
NAND_X1 U634 ( .A1(n600), .A2(n601), .A3(G11), .A4(n602), .ZN(G150) );
NOR_X1 U635 ( .A1(n603), .A2(n604), .ZN(n602) );
NOR_X1 U636 ( .A1(G29), .A2(n605), .ZN(n604) );
NOR_X1 U637 ( .A1(n606), .A2(n607), .ZN(n605) );
NAND_X1 U638 ( .A1(G28), .A2(n608), .A3(n609), .A4(n610), .ZN(w1095) );
XNOR_X1 U639 ( .A1(w1090), .A2(n500), .ZN(n610) );
INV_X1 U640 ( .A1(G2078), .ZN(n500) );
XNOR_X1 U641 ( .A1(w1092), .A2(n504), .ZN(n609) );
INV_X1 U642 ( .A1(G2084), .ZN(n504) );
XNOR_X1 U643 ( .A1(w1094), .A2(n508), .ZN(n608) );
INV_X1 U644 ( .A1(G2090), .ZN(n508) );
NAND_X1 U645 ( .A1(n611), .A2(n612), .A3(n613), .A4(n614), .ZN(w1101) );
XNOR_X1 U646 ( .A1(w1096), .A2(n551), .ZN(n614) );
XNOR_X1 U647 ( .A1(w1098), .A2(n441), .ZN(n613) );
XNOR_X1 U648 ( .A1(w1100), .A2(n434), .ZN(n612) );
INV_X1 U649 ( .A1(G2067), .ZN(n434) );
XOR_X1 U650 ( .A1(w1102), .A2(w1103), .ZN(n611) );
NOR_X1 U651 ( .A1(n615), .A2(n616), .ZN(n603) );
INV_X1 U652 ( .A1(G29), .ZN(n616) );
NOR_X1 U653 ( .A1(n617), .A2(n618), .A3(n515), .A4(n619), .ZN(w1105) );
XNOR_X1 U654 ( .A1(w1104), .A2(n510), .ZN(n619) );
NAND_X1 U655 ( .A1(n620), .A2(n621), .A3(n622), .A4(n623), .ZN(n510) );
NAND_X1 U656 ( .A1(G138), .A2(n573), .ZN(n623) );
NAND_X1 U657 ( .A1(G102), .A2(n574), .ZN(n622) );
NAND_X1 U658 ( .A1(G126), .A2(n575), .ZN(n621) );
NAND_X1 U659 ( .A1(G114), .A2(n576), .ZN(n620) );
NAND_X1 U660 ( .A1(n624), .A2(n625), .ZN(n515) );
NAND_X1 U661 ( .A1(G1991), .A2(n626), .ZN(n625) );
NAND_X1 U662 ( .A1(G1996), .A2(n627), .ZN(n624) );
NAND_X1 U663 ( .A1(n513), .A2(n556), .A3(n628), .ZN(n618) );
NAND_X1 U664 ( .A1(n440), .A2(n441), .ZN(n628) );
INV_X1 U665 ( .A1(G1996), .ZN(n441) );
INV_X1 U666 ( .A1(n627), .ZN(w1049) );
NAND_X1 U667 ( .A1(n629), .A2(n630), .A3(n631), .A4(n632), .ZN(n627) );
NAND_X1 U668 ( .A1(G141), .A2(n573), .ZN(n632) );
NAND_X1 U669 ( .A1(G105), .A2(n574), .ZN(n631) );
NAND_X1 U670 ( .A1(G129), .A2(n575), .ZN(n630) );
NAND_X1 U671 ( .A1(G117), .A2(n576), .ZN(n629) );
NAND_X1 U672 ( .A1(n633), .A2(n634), .A3(n635), .A4(n636), .ZN(n556) );
NAND_X1 U673 ( .A1(G135), .A2(n573), .ZN(n636) );
NAND_X1 U674 ( .A1(G99), .A2(n574), .ZN(n635) );
NAND_X1 U675 ( .A1(G123), .A2(n575), .ZN(n634) );
NAND_X1 U676 ( .A1(G111), .A2(n576), .ZN(n633) );
NAND_X1 U677 ( .A1(n567), .A2(n551), .ZN(n513) );
INV_X1 U678 ( .A1(G1991), .ZN(n551) );
INV_X1 U679 ( .A1(n626), .ZN(n567) );
NAND_X1 U680 ( .A1(n637), .A2(n638), .A3(n639), .A4(n640), .ZN(n626) );
NAND_X1 U681 ( .A1(G131), .A2(n573), .ZN(n640) );
NAND_X1 U682 ( .A1(G95), .A2(n574), .ZN(n639) );
NAND_X1 U683 ( .A1(G119), .A2(n575), .ZN(n638) );
NAND_X1 U684 ( .A1(G107), .A2(n576), .ZN(n637) );
NAND_X1 U685 ( .A1(n641), .A2(n642), .A3(n643), .A4(n644), .ZN(w1113) );
XNOR_X1 U686 ( .A1(G160), .A2(w1106), .ZN(n644) );
INV_X1 U687 ( .A1(n562), .ZN(G160) );
NAND_X1 U688 ( .A1(n645), .A2(n646), .A3(n647), .A4(n648), .ZN(w1043) );
NAND_X1 U689 ( .A1(G137), .A2(n573), .ZN(n648) );
NAND_X1 U690 ( .A1(G101), .A2(n574), .ZN(n647) );
NAND_X1 U691 ( .A1(G125), .A2(n575), .ZN(n646) );
NAND_X1 U692 ( .A1(G113), .A2(n576), .ZN(n645) );
XNOR_X1 U693 ( .A1(G162), .A2(w1108), .ZN(n643) );
AND_X1 U694 ( .A1(n649), .A2(n650), .A3(n651), .A4(n652), .ZN(G162) );
NAND_X1 U695 ( .A1(G136), .A2(n573), .ZN(n652) );
NAND_X1 U696 ( .A1(G100), .A2(n574), .ZN(n651) );
NAND_X1 U697 ( .A1(G124), .A2(n575), .ZN(n650) );
NAND_X1 U698 ( .A1(G112), .A2(n576), .ZN(n649) );
XOR_X1 U699 ( .A1(n563), .A2(w1110), .ZN(n642) );
NAND_X1 U700 ( .A1(n653), .A2(n654), .A3(n655), .A4(n656), .ZN(n563) );
NAND_X1 U701 ( .A1(G139), .A2(n573), .ZN(n656) );
NAND_X1 U702 ( .A1(G103), .A2(n574), .ZN(n655) );
NAND_X1 U703 ( .A1(G127), .A2(n575), .ZN(n654) );
NAND_X1 U704 ( .A1(G115), .A2(n576), .ZN(n653) );
XNOR_X1 U705 ( .A1(n437), .A2(w1112), .ZN(n641) );
INV_X1 U706 ( .A1(n566), .ZN(n437) );
NAND_X1 U707 ( .A1(n657), .A2(n658), .A3(n659), .A4(n660), .ZN(n566) );
NAND_X1 U708 ( .A1(G140), .A2(n573), .ZN(n660) );
NOR_X1 U709 ( .A1(G2104), .A2(G2105), .ZN(n573) );
NAND_X1 U710 ( .A1(G104), .A2(n574), .ZN(n659) );
NOR_X1 U711 ( .A1(n661), .A2(G2105), .ZN(n574) );
NAND_X1 U712 ( .A1(G128), .A2(n575), .ZN(n658) );
NOR_X1 U713 ( .A1(n662), .A2(G2104), .ZN(n575) );
NAND_X1 U714 ( .A1(G116), .A2(n576), .ZN(n657) );
NOR_X1 U715 ( .A1(n662), .A2(n661), .ZN(n576) );
INV_X1 U716 ( .A1(G2104), .ZN(n661) );
INV_X1 U717 ( .A1(G2105), .ZN(n662) );
NAND_X1 U718 ( .A1(G16), .A2(n663), .ZN(n601) );
NAND_X1 U719 ( .A1(n664), .A2(n665), .A3(n666), .A4(n667), .ZN(w1127) );
NOR_X1 U720 ( .A1(n668), .A2(n669), .A3(n670), .A4(n671), .ZN(w1117) );
XNOR_X1 U721 ( .A1(w1114), .A2(G286), .ZN(n671) );
NAND_X1 U722 ( .A1(n672), .A2(n673), .A3(n674), .A4(n675), .ZN(G286) );
NAND_X1 U723 ( .A1(G89), .A2(n676), .ZN(n675) );
NAND_X1 U724 ( .A1(G76), .A2(n677), .ZN(n674) );
NAND_X1 U725 ( .A1(G51), .A2(n678), .ZN(n673) );
NAND_X1 U726 ( .A1(G63), .A2(n679), .ZN(n672) );
NOR_X1 U727 ( .A1(G1976), .A2(G288), .ZN(n670) );
XNOR_X1 U728 ( .A1(w1116), .A2(n532), .ZN(n669) );
NAND_X1 U729 ( .A1(n491), .A2(n461), .A3(n680), .ZN(n668) );
NAND_X1 U730 ( .A1(G1348), .A2(n499), .ZN(n680) );
NAND_X1 U731 ( .A1(G1976), .A2(G288), .ZN(n461) );
NAND_X1 U732 ( .A1(n681), .A2(n682), .A3(n683), .A4(n684), .ZN(w1083) );
NAND_X1 U733 ( .A1(G49), .A2(n678), .ZN(n683) );
NAND_X1 U734 ( .A1(G87), .A2(n685), .ZN(n682) );
NAND_X1 U735 ( .A1(G74), .A2(G651), .ZN(n681) );
NAND_X1 U736 ( .A1(n686), .A2(n492), .ZN(n491) );
INV_X1 U737 ( .A1(G1348), .ZN(n492) );
NOR_X1 U738 ( .A1(n687), .A2(n688), .A3(n689), .ZN(w1123) );
XNOR_X1 U739 ( .A1(w1118), .A2(G290), .ZN(n689) );
NAND_X1 U740 ( .A1(n690), .A2(n691), .A3(n692), .A4(n693), .ZN(w1085) );
NAND_X1 U741 ( .A1(G85), .A2(n676), .ZN(n693) );
NAND_X1 U742 ( .A1(G72), .A2(n677), .ZN(n692) );
NAND_X1 U743 ( .A1(G47), .A2(n678), .ZN(n691) );
NAND_X1 U744 ( .A1(G60), .A2(n679), .ZN(n690) );
XNOR_X1 U745 ( .A1(w1120), .A2(G301), .ZN(n688) );
NAND_X1 U746 ( .A1(n694), .A2(n695), .A3(n696), .A4(n697), .ZN(G301) );
NAND_X1 U747 ( .A1(G90), .A2(n676), .ZN(n697) );
NAND_X1 U748 ( .A1(G77), .A2(n677), .ZN(n696) );
NAND_X1 U749 ( .A1(G52), .A2(n678), .ZN(n695) );
NAND_X1 U750 ( .A1(G64), .A2(n679), .ZN(n694) );
XNOR_X1 U751 ( .A1(w1122), .A2(G299), .ZN(n687) );
NAND_X1 U752 ( .A1(n698), .A2(n699), .A3(n700), .A4(n701), .ZN(G299) );
NAND_X1 U753 ( .A1(G91), .A2(n676), .ZN(n701) );
NAND_X1 U754 ( .A1(G78), .A2(n677), .ZN(n700) );
NAND_X1 U755 ( .A1(G53), .A2(n678), .ZN(n699) );
NAND_X1 U756 ( .A1(G65), .A2(n679), .ZN(n698) );
XNOR_X1 U757 ( .A1(G166), .A2(w1124), .ZN(n665) );
INV_X1 U758 ( .A1(G303), .ZN(G166) );
NAND_X1 U759 ( .A1(n702), .A2(n703), .A3(n704), .A4(n705), .ZN(G303) );
NAND_X1 U760 ( .A1(G88), .A2(n676), .ZN(n705) );
NAND_X1 U761 ( .A1(G75), .A2(n677), .ZN(n704) );
NAND_X1 U762 ( .A1(G50), .A2(n678), .ZN(n703) );
NAND_X1 U763 ( .A1(G62), .A2(n679), .ZN(n702) );
XOR_X1 U764 ( .A1(G305), .A2(w1126), .ZN(n664) );
NAND_X1 U765 ( .A1(n706), .A2(n707), .A3(n708), .A4(n709), .ZN(G305) );
NAND_X1 U766 ( .A1(G86), .A2(n676), .ZN(n709) );
NAND_X1 U767 ( .A1(G73), .A2(n677), .ZN(n708) );
NAND_X1 U768 ( .A1(G48), .A2(n678), .ZN(n707) );
NAND_X1 U769 ( .A1(G61), .A2(n679), .ZN(n706) );
NAND_X1 U770 ( .A1(n710), .A2(n711), .ZN(n600) );
INV_X1 U771 ( .A1(G16), .ZN(n711) );
NAND_X1 U772 ( .A1(n712), .A2(n713), .A3(n714), .A4(n715), .ZN(n710) );
NOR_X1 U773 ( .A1(n716), .A2(n717), .A3(n718), .A4(n719), .ZN(n715) );
XNOR_X1 U774 ( .A1(w1128), .A2(w1129), .ZN(n719) );
XNOR_X1 U775 ( .A1(w1130), .A2(w1131), .ZN(n718) );
XNOR_X1 U776 ( .A1(G1976), .A2(G23), .ZN(n717) );
XNOR_X1 U777 ( .A1(G1971), .A2(G22), .ZN(n716) );
NOR_X1 U778 ( .A1(n720), .A2(n721), .A3(n722), .ZN(n714) );
XNOR_X1 U779 ( .A1(G1341), .A2(G19), .ZN(n722) );
XNOR_X1 U780 ( .A1(G1956), .A2(G20), .ZN(n721) );
XNOR_X1 U781 ( .A1(G1348), .A2(G4), .ZN(n720) );
XNOR_X1 U782 ( .A1(G5), .A2(n501), .ZN(n713) );
INV_X1 U783 ( .A1(G1961), .ZN(n501) );
XNOR_X1 U784 ( .A1(G21), .A2(n505), .ZN(n712) );
INV_X1 U785 ( .A1(G1966), .ZN(n505) );
NAND_X1 U786 ( .A1(n686), .A2(n723), .ZN(G148) );
NAND_X1 U787 ( .A1(n526), .A2(n599), .ZN(n723) );
INV_X1 U788 ( .A1(n499), .ZN(n686) );
XNOR_X1 U789 ( .A1(n724), .A2(n522), .ZN(G145) );
NAND_X1 U790 ( .A1(n725), .A2(n726), .A3(n727), .A4(n728), .ZN(w1079) );
NAND_X1 U791 ( .A1(G93), .A2(n676), .ZN(n728) );
NAND_X1 U792 ( .A1(G80), .A2(n677), .ZN(n727) );
NAND_X1 U793 ( .A1(G55), .A2(n678), .ZN(n726) );
NAND_X1 U794 ( .A1(G67), .A2(n679), .ZN(n725) );
NAND_X1 U795 ( .A1(n486), .A2(n599), .A3(n729), .A4(n730), .ZN(n724) );
NAND_X1 U796 ( .A1(n731), .A2(n532), .ZN(n730) );
NAND_X1 U797 ( .A1(n493), .A2(n526), .ZN(n729) );
INV_X1 U798 ( .A1(n731), .ZN(n526) );
NOR_X1 U799 ( .A1(G559), .A2(n499), .ZN(n731) );
NOR_X1 U800 ( .A1(n532), .A2(n499), .ZN(n493) );
INV_X1 U801 ( .A1(G860), .ZN(n599) );
NAND_X1 U802 ( .A1(n532), .A2(n499), .ZN(n486) );
NAND_X1 U803 ( .A1(n732), .A2(n733), .A3(n734), .A4(n735), .ZN(n499) );
NAND_X1 U804 ( .A1(G92), .A2(n676), .ZN(n735) );
NAND_X1 U805 ( .A1(G79), .A2(n677), .ZN(n734) );
NAND_X1 U806 ( .A1(G54), .A2(n678), .ZN(n733) );
NAND_X1 U807 ( .A1(G66), .A2(n679), .ZN(n732) );
NAND_X1 U808 ( .A1(n736), .A2(n737), .A3(n738), .A4(n739), .ZN(n532) );
NAND_X1 U809 ( .A1(G81), .A2(n676), .ZN(n739) );
NOR_X1 U810 ( .A1(G543), .A2(G651), .ZN(n676) );
NAND_X1 U811 ( .A1(G68), .A2(n677), .ZN(n738) );
AND_X1 U812 ( .A1(G651), .A2(G543), .ZN(n677) );
NAND_X1 U813 ( .A1(G43), .A2(n678), .ZN(n737) );
NOR_X1 U814 ( .A1(n685), .A2(G651), .ZN(n678) );
NAND_X1 U815 ( .A1(G56), .A2(n679), .ZN(n736) );
INV_X1 U816 ( .A1(n684), .ZN(n679) );
NAND_X1 U817 ( .A1(G651), .A2(n685), .ZN(n684) );
INV_X1 U818 ( .A1(G543), .ZN(n685) );
XOR_X1 X1000 ( .A1(w1000), .A2(KEYINPUT0), .ZN(n520) );
XNOR_X1 X1001 ( .A1(w1001), .A2(KEYINPUT1), .ZN(n525) );
XOR_X1 X1002 ( .A1(w1002), .A2(KEYINPUT2), .ZN(n523) );
XNOR_X1 X1003 ( .A1(w1003), .A2(KEYINPUT3), .ZN(n527) );
XOR_X1 X1004 ( .A1(w1004), .A2(KEYINPUT4), .ZN(n536) );
XNOR_X1 X1005 ( .A1(w1005), .A2(KEYINPUT5), .ZN(n539) );
XOR_X1 X1006 ( .A1(w1006), .A2(KEYINPUT6), .ZN(G227) );
XNOR_X1 X1007 ( .A1(w1007), .A2(KEYINPUT7), .ZN(n541) );
XOR_X1 X1008 ( .A1(G2072), .A2(KEYINPUT8), .ZN(w1008) );
XNOR_X1 X1009 ( .A1(w1009), .A2(KEYINPUT9), .ZN(w1005) );
XOR_X1 X1010 ( .A1(G2078), .A2(KEYINPUT10), .ZN(w1010) );
XNOR_X1 X1011 ( .A1(w1011), .A2(KEYINPUT11), .ZN(w1009) );
XOR_X1 X1012 ( .A1(w1012), .A2(KEYINPUT12), .ZN(w1006) );
XNOR_X1 X1013 ( .A1(w1013), .A2(KEYINPUT13), .ZN(n543) );
XOR_X1 X1014 ( .A1(G2678), .A2(KEYINPUT14), .ZN(w1014) );
XNOR_X1 X1015 ( .A1(w1015), .A2(KEYINPUT15), .ZN(n538) );
XOR_X1 X1016 ( .A1(G2096), .A2(KEYINPUT16), .ZN(w1016) );
XNOR_X1 X1017 ( .A1(G2090), .A2(KEYINPUT17), .ZN(w1017) );
XOR_X1 X1018 ( .A1(w1018), .A2(KEYINPUT18), .ZN(w1004) );
XNOR_X1 X1019 ( .A1(w1019), .A2(KEYINPUT19), .ZN(n546) );
XOR_X1 X1020 ( .A1(G1986), .A2(KEYINPUT20), .ZN(w1020) );
XNOR_X1 X1021 ( .A1(G1981), .A2(KEYINPUT21), .ZN(w1021) );
XOR_X1 X1022 ( .A1(w1022), .A2(KEYINPUT22), .ZN(G229) );
XNOR_X1 X1023 ( .A1(w1023), .A2(KEYINPUT23), .ZN(n548) );
XOR_X1 X1024 ( .A1(w1024), .A2(KEYINPUT24), .ZN(n545) );
XNOR_X1 X1025 ( .A1(w1025), .A2(KEYINPUT25), .ZN(n550) );
XOR_X1 X1026 ( .A1(G1976), .A2(KEYINPUT26), .ZN(w1026) );
XNOR_X1 X1027 ( .A1(w1027), .A2(KEYINPUT27), .ZN(w1023) );
XOR_X1 X1028 ( .A1(G2474), .A2(KEYINPUT28), .ZN(w1028) );
XNOR_X1 X1029 ( .A1(w1029), .A2(KEYINPUT29), .ZN(w1027) );
XOR_X1 X1030 ( .A1(w1030), .A2(KEYINPUT30), .ZN(w1024) );
XNOR_X1 X1031 ( .A1(w1031), .A2(KEYINPUT31), .ZN(n553) );
XOR_X1 X1032 ( .A1(G1966), .A2(KEYINPUT32), .ZN(w1032) );
XNOR_X1 X1033 ( .A1(w1033), .A2(KEYINPUT33), .ZN(n547) );
XOR_X1 X1034 ( .A1(G1956), .A2(KEYINPUT34), .ZN(w1034) );
XNOR_X1 X1035 ( .A1(G1961), .A2(KEYINPUT35), .ZN(w1035) );
XOR_X1 X1036 ( .A1(w1036), .A2(KEYINPUT36), .ZN(n427) );
XNOR_X1 X1037 ( .A1(w1037), .A2(KEYINPUT37), .ZN(n557) );
XOR_X1 X1038 ( .A1(w1038), .A2(KEYINPUT38), .ZN(n554) );
XNOR_X1 X1039 ( .A1(w1039), .A2(KEYINPUT39), .ZN(n559) );
XOR_X1 X1040 ( .A1(w1040), .A2(KEYINPUT40), .ZN(w1037) );
XNOR_X1 X1041 ( .A1(w1041), .A2(KEYINPUT41), .ZN(n561) );
XOR_X1 X1042 ( .A1(w1042), .A2(KEYINPUT42), .ZN(w1039) );
XNOR_X1 X1043 ( .A1(w1043), .A2(KEYINPUT43), .ZN(n562) );
XOR_X1 X1044 ( .A1(w1044), .A2(KEYINPUT44), .ZN(w1042) );
XNOR_X1 X1045 ( .A1(w1045), .A2(KEYINPUT45), .ZN(G164) );
XOR_X1 X1046 ( .A1(w1046), .A2(KEYINPUT46), .ZN(w1040) );
XNOR_X1 X1047 ( .A1(w1047), .A2(KEYINPUT47), .ZN(n565) );
XOR_X1 X1048 ( .A1(w1048), .A2(KEYINPUT48), .ZN(n558) );
XNOR_X1 X1049 ( .A1(w1049), .A2(KEYINPUT49), .ZN(n440) );
XOR_X1 X1050 ( .A1(w1050), .A2(KEYINPUT50), .ZN(w1048) );
XNOR_X1 X1051 ( .A1(w1051), .A2(KEYINPUT51), .ZN(n568) );
XOR_X1 X1052 ( .A1(w1052), .A2(KEYINPUT52), .ZN(n425) );
XNOR_X1 X1053 ( .A1(w1053), .A2(KEYINPUT53), .ZN(n579) );
XOR_X1 X1054 ( .A1(G2430), .A2(KEYINPUT54), .ZN(w1054) );
XNOR_X1 X1055 ( .A1(G2427), .A2(KEYINPUT55), .ZN(w1055) );
XOR_X1 X1056 ( .A1(w1056), .A2(KEYINPUT56), .ZN(n577) );
XNOR_X1 X1057 ( .A1(w1057), .A2(KEYINPUT57), .ZN(n580) );
XOR_X1 X1058 ( .A1(w1058), .A2(KEYINPUT58), .ZN(n578) );
XNOR_X1 X1059 ( .A1(w1059), .A2(KEYINPUT59), .ZN(n582) );
XOR_X1 X1060 ( .A1(w1060), .A2(KEYINPUT60), .ZN(w1057) );
XNOR_X1 X1061 ( .A1(w1061), .A2(KEYINPUT61), .ZN(n584) );
XOR_X1 X1062 ( .A1(G2446), .A2(KEYINPUT62), .ZN(w1062) );
XNOR_X1 X1063 ( .A1(G2443), .A2(KEYINPUT63), .ZN(w1063) );
XOR_X1 X1064 ( .A1(G2454), .A2(KEYINPUT64), .ZN(w1064) );
XNOR_X1 X1065 ( .A1(G2451), .A2(KEYINPUT65), .ZN(w1065) );
XOR_X1 X1066 ( .A1(G1341), .A2(KEYINPUT66), .ZN(w1066) );
XNOR_X1 X1067 ( .A1(w1067), .A2(KEYINPUT67), .ZN(w1060) );
XOR_X1 X1068 ( .A1(G2438), .A2(KEYINPUT68), .ZN(w1068) );
XNOR_X1 X1069 ( .A1(G2435), .A2(KEYINPUT69), .ZN(w1069) );
XOR_X1 X1070 ( .A1(w1070), .A2(KEYINPUT70), .ZN(n426) );
XNOR_X1 X1071 ( .A1(w1071), .A2(KEYINPUT71), .ZN(n588) );
XOR_X1 X1072 ( .A1(w1072), .A2(KEYINPUT72), .ZN(n586) );
XNOR_X1 X1073 ( .A1(w1073), .A2(KEYINPUT73), .ZN(n589) );
XOR_X1 X1074 ( .A1(w1074), .A2(KEYINPUT74), .ZN(w1002) );
XNOR_X1 X1075 ( .A1(w1075), .A2(KEYINPUT75), .ZN(w1073) );
XOR_X1 X1076 ( .A1(w1076), .A2(KEYINPUT76), .ZN(n524) );
XNOR_X1 X1077 ( .A1(w1077), .A2(KEYINPUT77), .ZN(n481) );
XOR_X1 X1078 ( .A1(w1078), .A2(KEYINPUT78), .ZN(w1076) );
XNOR_X1 X1079 ( .A1(w1079), .A2(KEYINPUT79), .ZN(n522) );
XOR_X1 X1080 ( .A1(w1080), .A2(KEYINPUT80), .ZN(w1001) );
XNOR_X1 X1081 ( .A1(w1081), .A2(KEYINPUT81), .ZN(w1071) );
XOR_X1 X1082 ( .A1(w1082), .A2(KEYINPUT82), .ZN(w1003) );
XNOR_X1 X1083 ( .A1(w1083), .A2(KEYINPUT83), .ZN(G288) );
XOR_X1 X1084 ( .A1(w1084), .A2(KEYINPUT84), .ZN(w1082) );
XNOR_X1 X1085 ( .A1(w1085), .A2(KEYINPUT85), .ZN(G290) );
XOR_X1 X1086 ( .A1(w1086), .A2(KEYINPUT86), .ZN(w1072) );
XNOR_X1 X1087 ( .A1(w1087), .A2(KEYINPUT87), .ZN(G171) );
XOR_X1 X1088 ( .A1(G2096), .A2(KEYINPUT88), .ZN(w1088) );
XNOR_X1 X1089 ( .A1(w1089), .A2(KEYINPUT89), .ZN(G156) );
XOR_X1 X1090 ( .A1(G27), .A2(KEYINPUT90), .ZN(w1090) );
XNOR_X1 X1091 ( .A1(w1091), .A2(KEYINPUT91), .ZN(n607) );
XOR_X1 X1092 ( .A1(G34), .A2(KEYINPUT92), .ZN(w1092) );
XNOR_X1 X1093 ( .A1(w1093), .A2(KEYINPUT93), .ZN(w1091) );
XOR_X1 X1094 ( .A1(G35), .A2(KEYINPUT94), .ZN(w1094) );
XNOR_X1 X1095 ( .A1(w1095), .A2(KEYINPUT95), .ZN(w1093) );
XOR_X1 X1096 ( .A1(G25), .A2(KEYINPUT96), .ZN(w1096) );
XNOR_X1 X1097 ( .A1(w1097), .A2(KEYINPUT97), .ZN(n606) );
XOR_X1 X1098 ( .A1(G32), .A2(KEYINPUT98), .ZN(w1098) );
XNOR_X1 X1099 ( .A1(w1099), .A2(KEYINPUT99), .ZN(w1097) );
XOR_X1 X1100 ( .A1(G26), .A2(KEYINPUT100), .ZN(w1100) );
XNOR_X1 X1101 ( .A1(w1101), .A2(KEYINPUT101), .ZN(w1099) );
XOR_X1 X1102 ( .A1(G33), .A2(KEYINPUT102), .ZN(w1102) );
XNOR_X1 X1103 ( .A1(G2072), .A2(KEYINPUT103), .ZN(w1103) );
XOR_X1 X1104 ( .A1(G2078), .A2(KEYINPUT104), .ZN(w1104) );
XNOR_X1 X1105 ( .A1(w1105), .A2(KEYINPUT105), .ZN(n615) );
XOR_X1 X1106 ( .A1(G2084), .A2(KEYINPUT106), .ZN(w1106) );
XNOR_X1 X1107 ( .A1(w1107), .A2(KEYINPUT107), .ZN(n617) );
XOR_X1 X1108 ( .A1(G2090), .A2(KEYINPUT108), .ZN(w1108) );
XNOR_X1 X1109 ( .A1(w1109), .A2(KEYINPUT109), .ZN(w1107) );
XOR_X1 X1110 ( .A1(G2072), .A2(KEYINPUT110), .ZN(w1110) );
XNOR_X1 X1111 ( .A1(w1111), .A2(KEYINPUT111), .ZN(w1109) );
XOR_X1 X1112 ( .A1(G2067), .A2(KEYINPUT112), .ZN(w1112) );
XNOR_X1 X1113 ( .A1(w1113), .A2(KEYINPUT113), .ZN(w1111) );
XOR_X1 X1114 ( .A1(G1966), .A2(KEYINPUT114), .ZN(w1114) );
XNOR_X1 X1115 ( .A1(w1115), .A2(KEYINPUT115), .ZN(n667) );
XOR_X1 X1116 ( .A1(G1341), .A2(KEYINPUT116), .ZN(w1116) );
XNOR_X1 X1117 ( .A1(w1117), .A2(KEYINPUT117), .ZN(w1115) );
XOR_X1 X1118 ( .A1(G1986), .A2(KEYINPUT118), .ZN(w1118) );
XNOR_X1 X1119 ( .A1(w1119), .A2(KEYINPUT119), .ZN(n666) );
XOR_X1 X1120 ( .A1(G1961), .A2(KEYINPUT120), .ZN(w1120) );
XNOR_X1 X1121 ( .A1(w1121), .A2(KEYINPUT121), .ZN(w1119) );
XOR_X1 X1122 ( .A1(G1956), .A2(KEYINPUT122), .ZN(w1122) );
XNOR_X1 X1123 ( .A1(w1123), .A2(KEYINPUT123), .ZN(w1121) );
XOR_X1 X1124 ( .A1(G1971), .A2(KEYINPUT124), .ZN(w1124) );
XNOR_X1 X1125 ( .A1(w1125), .A2(KEYINPUT125), .ZN(n663) );
XOR_X1 X1126 ( .A1(G1981), .A2(KEYINPUT126), .ZN(w1126) );
XNOR_X1 X1127 ( .A1(w1127), .A2(KEYINPUT127), .ZN(w1125) );
XOR_X1 X1128 ( .A1(G1986), .A2(KEYINPUT128), .ZN(w1128) );
XNOR_X1 X1129 ( .A1(G24), .A2(KEYINPUT129), .ZN(w1129) );
XOR_X1 X1130 ( .A1(G1981), .A2(KEYINPUT130), .ZN(w1130) );
XNOR_X1 X1131 ( .A1(G6), .A2(KEYINPUT131), .ZN(w1131) );
