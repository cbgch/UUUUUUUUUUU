module c3540 ( G200,G213,G343,G2897,G326,G317,G294,G311,G303,G283,G329,G68,G97,G77,
G159,G50,G45,G322,G116,G58,G150,G143,G107,G330,G137,G87,G33,G20,
G132,G128,G125,G1,G13,G124,G190,G179,G238,G232,G226,G223,G222,G244,
G274,G41,G169,G264,G257,G270,G250,G1698,KEYINPUT0,KEYINPUT1,KEYINPUT2,KEYINPUT3,KEYINPUT4,KEYINPUT5,
KEYINPUT6,KEYINPUT7,KEYINPUT8,KEYINPUT9,KEYINPUT10,KEYINPUT11,KEYINPUT12,KEYINPUT13,KEYINPUT14,KEYINPUT15,KEYINPUT16,KEYINPUT17,KEYINPUT18,KEYINPUT19,
KEYINPUT20,KEYINPUT21,KEYINPUT22,KEYINPUT23,KEYINPUT24,KEYINPUT25,KEYINPUT26,KEYINPUT27,KEYINPUT28,KEYINPUT29,KEYINPUT30,KEYINPUT31,KEYINPUT32,KEYINPUT33,
KEYINPUT34,KEYINPUT35,KEYINPUT36,KEYINPUT37,KEYINPUT38,KEYINPUT39,KEYINPUT40,KEYINPUT41,KEYINPUT42,KEYINPUT43,KEYINPUT44,KEYINPUT45,KEYINPUT46,KEYINPUT47,
KEYINPUT48,KEYINPUT49,KEYINPUT50,KEYINPUT51,KEYINPUT52,KEYINPUT53,KEYINPUT54,KEYINPUT55,KEYINPUT56,KEYINPUT57,KEYINPUT58,KEYINPUT59,KEYINPUT60,KEYINPUT61,
KEYINPUT62,KEYINPUT63,KEYINPUT64,KEYINPUT65,KEYINPUT66,KEYINPUT67,KEYINPUT68,KEYINPUT69,KEYINPUT70,KEYINPUT71,KEYINPUT72,KEYINPUT73,KEYINPUT74,KEYINPUT75,
KEYINPUT76,KEYINPUT77,G409,G407,G405,G402,G396,G393,G390,G387,G399,G384,G381,G378,
G375,G372,G367,G369,G364,G361,G358,G355,G353,G351 );
input G200, G213, G343, G2897, G326,
 G317, G294, G311, G303, G283, G329, G68, G97, G77, G159, G50, G45, G322, G116,
 G58, G150, G143, G107, G330, G137, G87, G33, G20, G132, G128, G125, G1, G13,
 G124, G190, G179, G238, G232, G226, G223, G222, G244, G274, G41, G169, G264, G257,
 G270, G250, G1698, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
 KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
 KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
 KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
 KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65, KEYINPUT66,
 KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77;
output G409, G407, G405, G402, G396, G393, G390, G387, G399, G384, G381, G378, G375, G372,
 G367, G369, G364, G361, G358, G355, G353, G351;
NOR_X1 U1502 ( .A1(n2565), .A2(n2567), .A3(n2568), .ZN(n2208) );
NOR_X1 U1503 ( .A1(n2565), .A2(G200), .A3(n2566), .ZN(n2214) );
NOR_X1 U1504 ( .A1(n2568), .A2(n2565), .A3(n2566), .ZN(n2212) );
NAND_X1 U1505 ( .A1(n2172), .A2(G407), .A3(G213), .ZN(G409) );
OR_X1 U1506 ( .A1(G378), .A2(G343), .A3(G375), .ZN(n2172) );
NAND_X1 U1507 ( .A1(n2173), .A2(n2174), .A3(n2175), .A4(n2176), .ZN(G407) );
NOR_X1 U1508 ( .A1(G375), .A2(G384), .A3(G387), .A4(G396), .ZN(n2176) );
NOR_X1 U1509 ( .A1(G393), .A2(G390), .ZN(n2175) );
INV_X1 U1510 ( .A1(G381), .ZN(n2174) );
XOR_X1 U1511 ( .A1(n2177), .A2(n2178), .ZN(w1002) );
XOR_X1 U1512 ( .A1(n2179), .A2(n2180), .ZN(w1008) );
NOR_X1 U1513 ( .A1(n2181), .A2(n2173), .ZN(w1003) );
NAND_X1 U1514 ( .A1(n2182), .A2(n2183), .ZN(w1001) );
NAND_X1 U1515 ( .A1(G375), .A2(n2184), .ZN(n2183) );
NAND_X1 U1516 ( .A1(G2897), .A2(n2181), .ZN(n2182) );
INV_X1 U1517 ( .A1(n2184), .ZN(n2181) );
NAND_X1 U1518 ( .A1(G213), .A2(n2185), .ZN(n2184) );
XNOR_X1 U1519 ( .A1(n2186), .A2(G375), .ZN(w1006) );
XOR_X1 U1520 ( .A1(n2179), .A2(n2173), .ZN(w1009) );
INV_X1 U1521 ( .A1(G378), .ZN(w1007) );
XOR_X1 U1522 ( .A1(n2187), .A2(n2188), .ZN(w1014) );
XNOR_X1 U1523 ( .A1(G396), .A2(n2189), .ZN(w1012) );
XOR_X1 U1524 ( .A1(G384), .A2(G387), .ZN(w1011) );
XOR_X1 U1525 ( .A1(G381), .A2(n2190), .ZN(w1016) );
XOR_X1 U1526 ( .A1(G393), .A2(G390), .ZN(w1015) );
NAND_X1 U1527 ( .A1(n2191), .A2(n2192), .ZN(G396) );
NAND_X1 U1528 ( .A1(n2193), .A2(n2194), .ZN(w1019) );
XOR_X1 U1529 ( .A1(w1018), .A2(n2195), .ZN(n2193) );
NAND_X1 U1530 ( .A1(n2196), .A2(n2197), .A3(n2198), .A4(n2199), .ZN(n2191) );
NOR_X1 U1531 ( .A1(n2200), .A2(n2201), .ZN(n2198) );
NOR_X1 U1532 ( .A1(n2202), .A2(n2203), .A3(n2204), .A4(n2205), .ZN(n2201) );
NOR_X1 U1533 ( .A1(n2206), .A2(n2207), .ZN(n2205) );
AND_X1 U1534 ( .A1(n2208), .A2(G326), .ZN(n2204) );
NAND_X1 U1535 ( .A1(n2209), .A2(n2210), .A3(n2211), .ZN(n2203) );
NAND_X1 U1536 ( .A1(G317), .A2(n2212), .ZN(n2211) );
NAND_X1 U1537 ( .A1(G294), .A2(n2213), .ZN(n2210) );
NAND_X1 U1538 ( .A1(G311), .A2(n2214), .ZN(n2209) );
NAND_X1 U1539 ( .A1(n2215), .A2(n2216), .A3(n2217), .A4(n2218), .ZN(n2202) );
NAND_X1 U1540 ( .A1(G303), .A2(n2219), .ZN(n2218) );
NAND_X1 U1541 ( .A1(G283), .A2(n2220), .ZN(n2217) );
NAND_X1 U1542 ( .A1(G329), .A2(n2221), .ZN(n2216) );
NOR_X1 U1543 ( .A1(n2222), .A2(n2223), .A3(n2224), .A4(n2225), .ZN(n2200) );
NOR_X1 U1544 ( .A1(n2226), .A2(n2206), .ZN(n2225) );
NOR_X1 U1545 ( .A1(n2227), .A2(n2228), .ZN(n2224) );
NAND_X1 U1546 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(n2223) );
NAND_X1 U1547 ( .A1(n2212), .A2(G68), .ZN(n2231) );
NAND_X1 U1548 ( .A1(G97), .A2(n2213), .ZN(n2230) );
INV_X1 U1549 ( .A1(n2232), .ZN(n2213) );
NAND_X1 U1550 ( .A1(G77), .A2(n2214), .ZN(n2229) );
NAND_X1 U1551 ( .A1(n2233), .A2(n2234), .A3(n2235), .A4(n2236), .ZN(n2222) );
NAND_X1 U1552 ( .A1(n2221), .A2(G159), .ZN(n2234) );
NAND_X1 U1553 ( .A1(n2237), .A2(n2238), .ZN(n2197) );
NAND_X1 U1554 ( .A1(n2239), .A2(n2240), .A3(n2241), .ZN(n2238) );
NAND_X1 U1555 ( .A1(n2242), .A2(G355), .ZN(n2241) );
NAND_X1 U1556 ( .A1(n2243), .A2(n2244), .A3(n2245), .ZN(n2240) );
NAND_X1 U1557 ( .A1(n2246), .A2(n2247), .ZN(n2239) );
NAND_X1 U1558 ( .A1(n2248), .A2(n2249), .ZN(n2246) );
OR_X1 U1559 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
NAND_X1 U1560 ( .A1(n2252), .A2(n2251), .ZN(n2248) );
NAND_X1 U1561 ( .A1(n2253), .A2(n2254), .ZN(w1026) );
NAND_X1 U1562 ( .A1(n2255), .A2(n2256), .A3(n2257), .ZN(w1017) );
NAND_X1 U1563 ( .A1(n2199), .A2(n2258), .A3(n2259), .A4(n2260), .ZN(n2257) );
NAND_X1 U1564 ( .A1(n2237), .A2(n2261), .ZN(n2260) );
NAND_X1 U1565 ( .A1(n2262), .A2(n2263), .A3(n2264), .ZN(n2261) );
NAND_X1 U1566 ( .A1(n2242), .A2(n2265), .ZN(n2264) );
NAND_X1 U1567 ( .A1(n2243), .A2(n2266), .A3(n2245), .ZN(n2263) );
NAND_X1 U1568 ( .A1(n2247), .A2(n2267), .ZN(n2262) );
NAND_X1 U1569 ( .A1(n2268), .A2(n2269), .ZN(n2267) );
NAND_X1 U1570 ( .A1(n2270), .A2(n2251), .ZN(n2269) );
OR_X1 U1571 ( .A1(n2265), .A2(n2226), .A3(n2271), .A4(G50), .ZN(n2270) );
NAND_X1 U1572 ( .A1(n2272), .A2(G45), .ZN(w1054) );
NOR_X1 U1573 ( .A1(n2273), .A2(n2274), .ZN(n2259) );
NOR_X1 U1574 ( .A1(n2275), .A2(n2276), .A3(n2277), .A4(n2278), .ZN(n2274) );
NOR_X1 U1575 ( .A1(n2232), .A2(n2279), .ZN(n2278) );
NOR_X1 U1576 ( .A1(n2227), .A2(n2207), .ZN(n2277) );
INV_X1 U1577 ( .A1(G322), .ZN(n2207) );
NAND_X1 U1578 ( .A1(n2280), .A2(n2281), .A3(n2282), .ZN(n2276) );
NAND_X1 U1579 ( .A1(G311), .A2(n2212), .ZN(n2282) );
NAND_X1 U1580 ( .A1(G317), .A2(n2283), .ZN(n2281) );
NAND_X1 U1581 ( .A1(G303), .A2(n2214), .ZN(n2280) );
NAND_X1 U1582 ( .A1(n2215), .A2(n2284), .A3(n2285), .A4(n2286), .ZN(n2275) );
NAND_X1 U1583 ( .A1(G294), .A2(n2219), .ZN(n2286) );
NAND_X1 U1584 ( .A1(G116), .A2(n2220), .ZN(n2285) );
NAND_X1 U1585 ( .A1(G326), .A2(n2221), .ZN(n2284) );
NOR_X1 U1586 ( .A1(n2287), .A2(n2288), .A3(n2289), .A4(n2290), .ZN(n2273) );
NOR_X1 U1587 ( .A1(n2206), .A2(n2228), .ZN(n2289) );
NAND_X1 U1588 ( .A1(n2291), .A2(n2292), .A3(n2293), .ZN(n2288) );
NAND_X1 U1589 ( .A1(G58), .A2(n2212), .ZN(n2293) );
NAND_X1 U1590 ( .A1(G159), .A2(n2208), .ZN(n2292) );
NAND_X1 U1591 ( .A1(G68), .A2(n2214), .ZN(n2291) );
NAND_X1 U1592 ( .A1(n2233), .A2(n2294), .A3(n2295), .A4(n2296), .ZN(n2287) );
NAND_X1 U1593 ( .A1(G77), .A2(n2219), .ZN(n2296) );
NAND_X1 U1594 ( .A1(G150), .A2(n2221), .ZN(n2294) );
NAND_X1 U1595 ( .A1(n2254), .A2(n2297), .ZN(w1028) );
NAND_X1 U1596 ( .A1(n2298), .A2(n2299), .ZN(w1020) );
NAND_X1 U1597 ( .A1(n2300), .A2(n2301), .A3(n2302), .ZN(n2255) );
NAND_X1 U1598 ( .A1(n2303), .A2(n2304), .A3(n2305), .ZN(G390) );
NAND_X1 U1599 ( .A1(n2306), .A2(n2299), .ZN(w1022) );
NAND_X1 U1600 ( .A1(n2307), .A2(n2308), .ZN(n2299) );
NAND_X1 U1601 ( .A1(n2300), .A2(n2309), .ZN(n2308) );
NAND_X1 U1602 ( .A1(n2310), .A2(n2311), .A3(n2199), .A4(n2312), .ZN(n2304) );
NOR_X1 U1603 ( .A1(n2313), .A2(n2242), .A3(n2314), .ZN(n2312) );
NOR_X1 U1604 ( .A1(n2315), .A2(n2316), .A3(n2317), .A4(n2318), .ZN(n2314) );
NOR_X1 U1605 ( .A1(n2319), .A2(n2206), .ZN(n2317) );
NAND_X1 U1606 ( .A1(n2320), .A2(n2321), .A3(n2322), .ZN(n2316) );
NAND_X1 U1607 ( .A1(G50), .A2(n2212), .ZN(n2322) );
NAND_X1 U1608 ( .A1(G150), .A2(n2208), .ZN(n2321) );
NAND_X1 U1609 ( .A1(G58), .A2(n2214), .ZN(n2320) );
NAND_X1 U1610 ( .A1(n2233), .A2(n2323), .A3(n2324), .A4(n2325), .ZN(n2315) );
NAND_X1 U1611 ( .A1(n2219), .A2(G68), .ZN(n2325) );
NAND_X1 U1612 ( .A1(G143), .A2(n2221), .ZN(n2323) );
NOR_X1 U1613 ( .A1(n2326), .A2(n2327), .A3(n2328), .A4(n2329), .ZN(n2313) );
NOR_X1 U1614 ( .A1(n2232), .A2(n2244), .ZN(n2329) );
AND_X1 U1615 ( .A1(n2208), .A2(G317), .ZN(n2328) );
NAND_X1 U1616 ( .A1(n2330), .A2(n2331), .A3(n2332), .ZN(n2327) );
NAND_X1 U1617 ( .A1(G303), .A2(n2212), .ZN(n2332) );
NAND_X1 U1618 ( .A1(G311), .A2(n2283), .ZN(n2331) );
NAND_X1 U1619 ( .A1(G294), .A2(n2214), .ZN(n2330) );
NAND_X1 U1620 ( .A1(n2215), .A2(n2333), .A3(n2235), .A4(n2334), .ZN(n2326) );
NAND_X1 U1621 ( .A1(G283), .A2(n2219), .ZN(n2334) );
NAND_X1 U1622 ( .A1(G107), .A2(n2220), .ZN(n2235) );
NAND_X1 U1623 ( .A1(G322), .A2(n2221), .ZN(n2333) );
NAND_X1 U1624 ( .A1(n2335), .A2(n2336), .A3(n2237), .ZN(n2311) );
NAND_X1 U1625 ( .A1(G97), .A2(n2245), .ZN(n2336) );
OR_X1 U1626 ( .A1(n2245), .A2(n2337), .ZN(w1068) );
NAND_X1 U1627 ( .A1(n2338), .A2(n2254), .ZN(w1030) );
NAND_X1 U1628 ( .A1(n2339), .A2(n2340), .A3(n2300), .ZN(n2303) );
NAND_X1 U1629 ( .A1(n2298), .A2(n2341), .ZN(w1021) );
NAND_X1 U1630 ( .A1(n2301), .A2(n2342), .ZN(n2341) );
NAND_X1 U1631 ( .A1(n2302), .A2(n2342), .ZN(n2339) );
INV_X1 U1632 ( .A1(n2306), .ZN(w1023) );
INV_X1 U1633 ( .A1(n2298), .ZN(n2302) );
NAND_X1 U1634 ( .A1(n2343), .A2(n2344), .ZN(w1013) );
NAND_X1 U1635 ( .A1(n2345), .A2(n2346), .A3(n2194), .ZN(w1024) );
NAND_X1 U1636 ( .A1(n2307), .A2(n2347), .A3(n2301), .ZN(n2346) );
NAND_X1 U1637 ( .A1(n2306), .A2(n2298), .ZN(n2347) );
XOR_X1 U1638 ( .A1(n2348), .A2(n2349), .ZN(n2298) );
XOR_X1 U1639 ( .A1(G399), .A2(n2350), .ZN(n2306) );
XNOR_X1 U1640 ( .A1(n2351), .A2(n2352), .ZN(w1032) );
NAND_X1 U1641 ( .A1(n2353), .A2(n2354), .ZN(w1025) );
NAND_X1 U1642 ( .A1(n2350), .A2(G399), .ZN(n2354) );
NAND_X1 U1643 ( .A1(n2355), .A2(n2356), .ZN(G399) );
NAND_X1 U1644 ( .A1(n2349), .A2(n2348), .ZN(n2356) );
NAND_X1 U1645 ( .A1(n2357), .A2(n2358), .ZN(n2348) );
NAND_X1 U1646 ( .A1(G330), .A2(n2195), .ZN(n2358) );
INV_X1 U1647 ( .A1(n2253), .ZN(w1027) );
XOR_X1 U1648 ( .A1(n2359), .A2(n2360), .ZN(n2253) );
NOR_X1 U1649 ( .A1(n2361), .A2(n2362), .ZN(n2360) );
OR_X1 U1650 ( .A1(n2363), .A2(n2364), .ZN(n2357) );
INV_X1 U1651 ( .A1(n2297), .ZN(w1029) );
XOR_X1 U1652 ( .A1(n2365), .A2(n2366), .ZN(n2297) );
NOR_X1 U1653 ( .A1(n2367), .A2(n2362), .ZN(n2366) );
OR_X1 U1654 ( .A1(n2368), .A2(n2364), .ZN(n2355) );
INV_X1 U1655 ( .A1(n2338), .ZN(w1031) );
XOR_X1 U1656 ( .A1(n2369), .A2(n2370), .ZN(n2338) );
NOR_X1 U1657 ( .A1(n2371), .A2(n2362), .ZN(n2370) );
OR_X1 U1658 ( .A1(n2372), .A2(n2364), .ZN(n2353) );
NAND_X1 U1659 ( .A1(n2373), .A2(n2374), .A3(n2375), .A4(n2199), .ZN(n2343) );
NOR_X1 U1660 ( .A1(n2376), .A2(n2242), .A3(n2377), .ZN(n2375) );
NOR_X1 U1661 ( .A1(n2378), .A2(n2379), .A3(n2380), .A4(n2381), .ZN(n2377) );
NOR_X1 U1662 ( .A1(n2232), .A2(n2266), .ZN(n2381) );
NOR_X1 U1663 ( .A1(n2206), .A2(n2382), .ZN(n2380) );
NAND_X1 U1664 ( .A1(n2383), .A2(n2384), .A3(n2385), .ZN(n2379) );
NAND_X1 U1665 ( .A1(G294), .A2(n2212), .ZN(n2385) );
NAND_X1 U1666 ( .A1(G311), .A2(n2208), .ZN(n2384) );
NAND_X1 U1667 ( .A1(G283), .A2(n2214), .ZN(n2383) );
NAND_X1 U1668 ( .A1(n2215), .A2(n2386), .A3(n2295), .A4(n2387), .ZN(n2378) );
NAND_X1 U1669 ( .A1(G116), .A2(n2219), .ZN(n2387) );
NAND_X1 U1670 ( .A1(G97), .A2(n2220), .ZN(n2295) );
NAND_X1 U1671 ( .A1(G317), .A2(n2221), .ZN(n2386) );
INV_X1 U1672 ( .A1(n2243), .ZN(n2242) );
NAND_X1 U1673 ( .A1(n2388), .A2(n2389), .ZN(n2243) );
NOR_X1 U1674 ( .A1(n2390), .A2(n2391), .A3(n2392), .A4(n2393), .ZN(n2376) );
NOR_X1 U1675 ( .A1(n2206), .A2(n2394), .ZN(n2392) );
NAND_X1 U1676 ( .A1(n2395), .A2(n2396), .A3(n2397), .ZN(n2391) );
NAND_X1 U1677 ( .A1(n2212), .A2(G159), .ZN(n2397) );
NAND_X1 U1678 ( .A1(G143), .A2(n2208), .ZN(n2396) );
NAND_X1 U1679 ( .A1(G50), .A2(n2214), .ZN(n2395) );
NAND_X1 U1680 ( .A1(n2233), .A2(n2398), .A3(n2399), .A4(n2400), .ZN(n2390) );
NAND_X1 U1681 ( .A1(n2219), .A2(G58), .ZN(n2400) );
NAND_X1 U1682 ( .A1(G137), .A2(n2221), .ZN(n2398) );
NAND_X1 U1683 ( .A1(n2401), .A2(n2402), .A3(n2237), .ZN(n2374) );
NOR_X1 U1684 ( .A1(n2403), .A2(n2254), .ZN(n2237) );
NAND_X1 U1685 ( .A1(G87), .A2(n2245), .ZN(n2402) );
NAND_X1 U1686 ( .A1(n2247), .A2(n2404), .ZN(w1060) );
INV_X1 U1687 ( .A1(n2245), .ZN(n2247) );
NAND_X1 U1688 ( .A1(G33), .A2(n2388), .ZN(n2245) );
NAND_X1 U1689 ( .A1(n2352), .A2(n2254), .ZN(w1033) );
NOR_X1 U1690 ( .A1(n2405), .A2(G20), .ZN(n2254) );
XNOR_X1 U1691 ( .A1(n2406), .A2(n2407), .ZN(n2352) );
NOR_X1 U1692 ( .A1(n2408), .A2(n2362), .ZN(n2407) );
NAND_X1 U1693 ( .A1(n2409), .A2(n2410), .ZN(G384) );
NAND_X1 U1694 ( .A1(n2411), .A2(n2194), .ZN(w1034) );
XOR_X1 U1695 ( .A1(n2301), .A2(n2412), .ZN(w1048) );
INV_X1 U1696 ( .A1(n2309), .ZN(w1035) );
NAND_X1 U1697 ( .A1(n2413), .A2(n2414), .A3(n2415), .A4(n2199), .ZN(n2409) );
NOR_X1 U1698 ( .A1(n2416), .A2(n2417), .ZN(n2415) );
NOR_X1 U1699 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(n2417) );
NOR_X1 U1700 ( .A1(n2226), .A2(n2232), .ZN(n2421) );
NOR_X1 U1701 ( .A1(n2206), .A2(n2422), .ZN(n2420) );
NAND_X1 U1702 ( .A1(n2423), .A2(n2424), .A3(n2425), .ZN(n2419) );
NAND_X1 U1703 ( .A1(G150), .A2(n2212), .ZN(n2425) );
NAND_X1 U1704 ( .A1(G137), .A2(n2208), .ZN(n2424) );
NAND_X1 U1705 ( .A1(n2214), .A2(G159), .ZN(n2423) );
NAND_X1 U1706 ( .A1(n2233), .A2(n2426), .A3(n2427), .A4(n2428), .ZN(n2418) );
NAND_X1 U1707 ( .A1(n2219), .A2(G50), .ZN(n2428) );
NAND_X1 U1708 ( .A1(G132), .A2(n2221), .ZN(n2426) );
NOR_X1 U1709 ( .A1(n2429), .A2(n2430), .A3(n2431), .A4(n2432), .ZN(n2416) );
NOR_X1 U1710 ( .A1(n2232), .A2(n2433), .ZN(n2432) );
NOR_X1 U1711 ( .A1(n2227), .A2(n2382), .ZN(n2431) );
INV_X1 U1712 ( .A1(G303), .ZN(n2382) );
NAND_X1 U1713 ( .A1(n2434), .A2(n2435), .A3(n2436), .ZN(n2430) );
NAND_X1 U1714 ( .A1(G283), .A2(n2212), .ZN(n2436) );
NAND_X1 U1715 ( .A1(G294), .A2(n2283), .ZN(n2435) );
NAND_X1 U1716 ( .A1(G116), .A2(n2214), .ZN(n2434) );
NAND_X1 U1717 ( .A1(n2215), .A2(n2437), .A3(n2324), .A4(n2438), .ZN(n2429) );
NAND_X1 U1718 ( .A1(G107), .A2(n2219), .ZN(n2438) );
NAND_X1 U1719 ( .A1(n2220), .A2(G87), .ZN(n2324) );
NAND_X1 U1720 ( .A1(G311), .A2(n2221), .ZN(n2437) );
NAND_X1 U1721 ( .A1(n2439), .A2(n2440), .ZN(n2414) );
NAND_X1 U1722 ( .A1(n2412), .A2(n2441), .ZN(w1049) );
NAND_X1 U1723 ( .A1(n2442), .A2(n2443), .A3(n2444), .ZN(G381) );
NAND_X1 U1724 ( .A1(n2199), .A2(n2445), .A3(n2446), .A4(n2447), .ZN(n2444) );
NAND_X1 U1725 ( .A1(n2439), .A2(n2448), .ZN(n2447) );
NOR_X1 U1726 ( .A1(n2449), .A2(n2450), .ZN(n2446) );
NOR_X1 U1727 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2450) );
NOR_X1 U1728 ( .A1(n2228), .A2(n2232), .ZN(n2454) );
NOR_X1 U1729 ( .A1(n2206), .A2(n2455), .ZN(n2453) );
NAND_X1 U1730 ( .A1(n2456), .A2(n2457), .A3(n2458), .ZN(n2452) );
NAND_X1 U1731 ( .A1(G143), .A2(n2212), .ZN(n2458) );
NAND_X1 U1732 ( .A1(G132), .A2(n2208), .ZN(n2457) );
NAND_X1 U1733 ( .A1(G150), .A2(n2214), .ZN(n2456) );
NAND_X1 U1734 ( .A1(n2233), .A2(n2459), .A3(n2460), .A4(n2461), .ZN(n2451) );
NAND_X1 U1735 ( .A1(n2219), .A2(G159), .ZN(n2461) );
NAND_X1 U1736 ( .A1(n2220), .A2(G58), .ZN(n2460) );
NAND_X1 U1737 ( .A1(G128), .A2(n2221), .ZN(n2459) );
NOR_X1 U1738 ( .A1(n2462), .A2(n2463), .A3(n2464), .A4(n2290), .ZN(n2449) );
NOR_X1 U1739 ( .A1(n2232), .A2(n2465), .ZN(n2290) );
AND_X1 U1740 ( .A1(n2208), .A2(G294), .ZN(n2464) );
NAND_X1 U1741 ( .A1(n2466), .A2(n2467), .A3(n2468), .ZN(n2463) );
NAND_X1 U1742 ( .A1(G116), .A2(n2212), .ZN(n2468) );
NAND_X1 U1743 ( .A1(G283), .A2(n2283), .ZN(n2467) );
NAND_X1 U1744 ( .A1(G107), .A2(n2214), .ZN(n2466) );
NAND_X1 U1745 ( .A1(n2215), .A2(n2469), .A3(n2399), .A4(n2470), .ZN(n2462) );
NAND_X1 U1746 ( .A1(G97), .A2(n2219), .ZN(n2470) );
NAND_X1 U1747 ( .A1(n2220), .A2(G77), .ZN(n2399) );
NAND_X1 U1748 ( .A1(G303), .A2(n2221), .ZN(n2469) );
NAND_X1 U1749 ( .A1(n2471), .A2(n2441), .ZN(w1050) );
NAND_X1 U1750 ( .A1(n2472), .A2(n2473), .ZN(n2443) );
NAND_X1 U1751 ( .A1(n2474), .A2(n2300), .A3(n2475), .ZN(n2442) );
NAND_X1 U1752 ( .A1(n2476), .A2(n2477), .A3(n2478), .ZN(G378) );
NAND_X1 U1753 ( .A1(n2479), .A2(n2473), .ZN(w1036) );
NAND_X1 U1754 ( .A1(n2307), .A2(n2480), .ZN(n2473) );
NAND_X1 U1755 ( .A1(n2300), .A2(n2481), .ZN(n2480) );
NAND_X1 U1756 ( .A1(n2199), .A2(n2482), .A3(n2483), .A4(n2484), .ZN(n2477) );
NAND_X1 U1757 ( .A1(n2439), .A2(n2226), .ZN(n2484) );
NOR_X1 U1758 ( .A1(n2403), .A2(n2441), .ZN(n2439) );
NOR_X1 U1759 ( .A1(n2485), .A2(n2486), .ZN(n2483) );
NOR_X1 U1760 ( .A1(n2487), .A2(n2488), .A3(n2489), .A4(n2490), .ZN(n2486) );
NOR_X1 U1761 ( .A1(n2319), .A2(n2232), .ZN(n2490) );
AND_X1 U1762 ( .A1(n2283), .A2(G132), .ZN(n2489) );
NAND_X1 U1763 ( .A1(n2491), .A2(n2492), .A3(n2493), .ZN(n2488) );
NAND_X1 U1764 ( .A1(G137), .A2(n2212), .ZN(n2493) );
NAND_X1 U1765 ( .A1(G128), .A2(n2208), .ZN(n2492) );
NAND_X1 U1766 ( .A1(G143), .A2(n2214), .ZN(n2491) );
NAND_X1 U1767 ( .A1(n2233), .A2(n2494), .A3(n2495), .A4(n2496), .ZN(n2487) );
NAND_X1 U1768 ( .A1(G150), .A2(n2219), .ZN(n2496) );
NAND_X1 U1769 ( .A1(n2220), .A2(G50), .ZN(n2495) );
NAND_X1 U1770 ( .A1(G125), .A2(n2221), .ZN(n2494) );
INV_X1 U1771 ( .A1(n2497), .ZN(n2233) );
NOR_X1 U1772 ( .A1(n2498), .A2(n2499), .A3(n2500), .A4(n2318), .ZN(n2485) );
NOR_X1 U1773 ( .A1(n2232), .A2(n2440), .ZN(n2318) );
NOR_X1 U1774 ( .A1(n2227), .A2(n2279), .ZN(n2500) );
INV_X1 U1775 ( .A1(G283), .ZN(n2279) );
INV_X1 U1776 ( .A1(n2208), .ZN(n2227) );
NAND_X1 U1777 ( .A1(n2501), .A2(n2502), .A3(n2503), .ZN(n2499) );
NAND_X1 U1778 ( .A1(G107), .A2(n2212), .ZN(n2503) );
NAND_X1 U1779 ( .A1(G116), .A2(n2283), .ZN(n2502) );
NAND_X1 U1780 ( .A1(G97), .A2(n2214), .ZN(n2501) );
NAND_X1 U1781 ( .A1(n2215), .A2(n2504), .A3(n2427), .A4(n2236), .ZN(n2498) );
NAND_X1 U1782 ( .A1(n2219), .A2(G87), .ZN(n2236) );
INV_X1 U1783 ( .A1(n2505), .ZN(n2219) );
NAND_X1 U1784 ( .A1(n2220), .A2(G68), .ZN(n2427) );
INV_X1 U1785 ( .A1(n2506), .ZN(n2220) );
NAND_X1 U1786 ( .A1(G294), .A2(n2221), .ZN(n2504) );
INV_X1 U1787 ( .A1(n2507), .ZN(n2215) );
NAND_X1 U1788 ( .A1(n2508), .A2(n2441), .ZN(w1046) );
INV_X1 U1789 ( .A1(n2405), .ZN(n2441) );
NAND_X1 U1790 ( .A1(n2509), .A2(n2510), .A3(n2300), .ZN(n2476) );
NAND_X1 U1791 ( .A1(n2472), .A2(n2511), .ZN(n2510) );
NAND_X1 U1792 ( .A1(n2474), .A2(n2512), .ZN(n2511) );
NAND_X1 U1793 ( .A1(n2512), .A2(n2475), .ZN(n2509) );
INV_X1 U1794 ( .A1(n2479), .ZN(w1037) );
NAND_X1 U1795 ( .A1(n2513), .A2(n2514), .ZN(w1005) );
NAND_X1 U1796 ( .A1(n2515), .A2(n2516), .A3(n2194), .ZN(w1038) );
INV_X1 U1797 ( .A1(n2199), .ZN(n2194) );
NAND_X1 U1798 ( .A1(n2307), .A2(n2517), .A3(n2474), .ZN(n2516) );
INV_X1 U1799 ( .A1(n2481), .ZN(n2474) );
NAND_X1 U1800 ( .A1(n2518), .A2(n2519), .ZN(n2481) );
OR_X1 U1801 ( .A1(n2520), .A2(n2521), .ZN(n2519) );
NAND_X1 U1802 ( .A1(n2479), .A2(n2472), .ZN(n2517) );
INV_X1 U1803 ( .A1(n2475), .ZN(n2472) );
NAND_X1 U1804 ( .A1(n2522), .A2(n2523), .ZN(n2475) );
NAND_X1 U1805 ( .A1(n2471), .A2(n2524), .ZN(w1051) );
NAND_X1 U1806 ( .A1(n2525), .A2(n2526), .ZN(n2524) );
NAND_X1 U1807 ( .A1(n2527), .A2(n2521), .ZN(n2526) );
NAND_X1 U1808 ( .A1(n2412), .A2(n2528), .ZN(n2525) );
XOR_X1 U1809 ( .A1(n2529), .A2(n2530), .ZN(n2479) );
NAND_X1 U1810 ( .A1(n2522), .A2(n2531), .ZN(n2529) );
NOR_X1 U1811 ( .A1(n2532), .A2(n2533), .ZN(n2522) );
INV_X1 U1812 ( .A1(n2534), .ZN(n2307) );
XOR_X1 U1813 ( .A1(n2535), .A2(n2536), .ZN(w1040) );
NAND_X1 U1814 ( .A1(n2537), .A2(n2538), .ZN(w1039) );
NAND_X1 U1815 ( .A1(n2539), .A2(n2540), .A3(n2541), .A4(n2199), .ZN(n2513) );
NOR_X1 U1816 ( .A1(n2534), .A2(n2300), .ZN(n2199) );
NAND_X1 U1817 ( .A1(G1), .A2(n2542), .ZN(n2534) );
NAND_X1 U1818 ( .A1(G13), .A2(n2543), .A3(G45), .ZN(n2542) );
NAND_X1 U1819 ( .A1(n2544), .A2(n2545), .ZN(n2541) );
NAND_X1 U1820 ( .A1(n2546), .A2(n2547), .ZN(n2544) );
NAND_X1 U1821 ( .A1(n2548), .A2(n2549), .A3(n2550), .A4(n2551), .ZN(n2547) );
NOR_X1 U1822 ( .A1(n2552), .A2(n2553), .A3(n2554), .A4(n2507), .ZN(n2551) );
NAND_X1 U1823 ( .A1(G33), .A2(n2403), .ZN(n2507) );
AND_X1 U1824 ( .A1(n2212), .A2(G97), .ZN(n2554) );
NOR_X1 U1825 ( .A1(n2505), .A2(n2440), .ZN(n2553) );
NOR_X1 U1826 ( .A1(n2206), .A2(n2266), .ZN(n2552) );
INV_X1 U1827 ( .A1(n2283), .ZN(n2206) );
NOR_X1 U1828 ( .A1(n2555), .A2(n2556), .A3(n2393), .ZN(n2550) );
NOR_X1 U1829 ( .A1(n2448), .A2(n2232), .ZN(n2393) );
NOR_X1 U1830 ( .A1(n2557), .A2(n2465), .ZN(n2556) );
NOR_X1 U1831 ( .A1(n2226), .A2(n2506), .ZN(n2555) );
NAND_X1 U1832 ( .A1(G283), .A2(n2221), .ZN(n2549) );
NAND_X1 U1833 ( .A1(G116), .A2(n2208), .ZN(n2548) );
NAND_X1 U1834 ( .A1(n2558), .A2(n2559), .A3(n2560), .A4(n2561), .ZN(n2546) );
NOR_X1 U1835 ( .A1(n2562), .A2(n2563), .A3(n2564), .A4(n2497), .ZN(n2561) );
NAND_X1 U1836 ( .A1(n2403), .A2(n2389), .ZN(n2497) );
NOR_X1 U1837 ( .A1(n2557), .A2(n2455), .ZN(n2564) );
INV_X1 U1838 ( .A1(G137), .ZN(n2455) );
INV_X1 U1839 ( .A1(n2214), .ZN(n2557) );
AND_X1 U1840 ( .A1(n2283), .A2(G128), .ZN(n2563) );
NOR_X1 U1841 ( .A1(n2567), .A2(G200), .A3(n2565), .ZN(n2283) );
AND_X1 U1842 ( .A1(n2208), .A2(G125), .ZN(n2562) );
NOR_X1 U1843 ( .A1(n2569), .A2(n2570), .A3(n2571), .ZN(n2560) );
NOR_X1 U1844 ( .A1(n2505), .A2(n2422), .ZN(n2571) );
INV_X1 U1845 ( .A1(G143), .ZN(n2422) );
NAND_X1 U1846 ( .A1(G200), .A2(G20), .A3(n2565), .A4(n2566), .ZN(n2505) );
NOR_X1 U1847 ( .A1(n2232), .A2(n2394), .ZN(n2570) );
NAND_X1 U1848 ( .A1(n2572), .A2(n2566), .ZN(n2232) );
NOR_X1 U1849 ( .A1(n2319), .A2(n2506), .ZN(n2569) );
NAND_X1 U1850 ( .A1(G200), .A2(n2565), .A3(n2567), .ZN(n2506) );
NAND_X1 U1851 ( .A1(G124), .A2(n2221), .ZN(n2559) );
AND_X1 U1852 ( .A1(n2572), .A2(n2567), .ZN(n2221) );
AND_X1 U1853 ( .A1(n2565), .A2(n2573), .ZN(n2572) );
NAND_X1 U1854 ( .A1(G200), .A2(G20), .ZN(n2573) );
NAND_X1 U1855 ( .A1(G132), .A2(n2212), .ZN(n2558) );
INV_X1 U1856 ( .A1(n2567), .ZN(n2566) );
NOR_X1 U1857 ( .A1(n2543), .A2(G190), .ZN(n2567) );
NAND_X1 U1858 ( .A1(G179), .A2(G20), .ZN(n2565) );
INV_X1 U1859 ( .A1(G200), .ZN(n2568) );
NAND_X1 U1860 ( .A1(n2574), .A2(n2228), .A3(n2405), .ZN(n2540) );
NAND_X1 U1861 ( .A1(n2403), .A2(n2545), .ZN(n2574) );
AND_X1 U1862 ( .A1(G13), .A2(n2575), .ZN(n2403) );
NAND_X1 U1863 ( .A1(G20), .A2(n2576), .ZN(n2575) );
OR_X1 U1864 ( .A1(n2536), .A2(n2405), .ZN(w1041) );
XNOR_X1 U1865 ( .A1(n2577), .A2(n2578), .ZN(n2536) );
NOR_X1 U1866 ( .A1(n2579), .A2(n2580), .ZN(n2578) );
NOR_X1 U1867 ( .A1(n2520), .A2(n2581), .ZN(G372) );
NAND_X1 U1868 ( .A1(n2582), .A2(n2583), .A3(n2584), .ZN(G367) );
NAND_X1 U1869 ( .A1(n2585), .A2(n2586), .A3(G1), .ZN(n2584) );
NAND_X1 U1870 ( .A1(n2587), .A2(n2588), .A3(n2589), .ZN(n2585) );
NAND_X1 U1871 ( .A1(G68), .A2(n2228), .ZN(n2589) );
NAND_X1 U1872 ( .A1(G50), .A2(n2448), .A3(G77), .A4(G58), .ZN(n2588) );
NAND_X1 U1873 ( .A1(n2271), .A2(n2226), .ZN(n2587) );
NAND_X1 U1874 ( .A1(n2590), .A2(n2591), .A3(n2592), .ZN(w1042) );
NAND_X1 U1875 ( .A1(G1), .A2(n2586), .ZN(n2591) );
XOR_X1 U1876 ( .A1(n2593), .A2(n2594), .ZN(w1044) );
XNOR_X1 U1877 ( .A1(n2537), .A2(n2518), .ZN(w1043) );
NAND_X1 U1878 ( .A1(G369), .A2(n2595), .ZN(w1045) );
NAND_X1 U1879 ( .A1(n2596), .A2(n2364), .ZN(n2595) );
NAND_X1 U1880 ( .A1(n2596), .A2(n2597), .ZN(G369) );
NAND_X1 U1881 ( .A1(n2598), .A2(n2599), .ZN(n2597) );
AND_X1 U1882 ( .A1(n2600), .A2(n2601), .ZN(n2596) );
NAND_X1 U1883 ( .A1(n2602), .A2(n2603), .ZN(n2600) );
NAND_X1 U1884 ( .A1(n2604), .A2(n2605), .ZN(n2603) );
NAND_X1 U1885 ( .A1(n2606), .A2(n2607), .ZN(n2604) );
NAND_X1 U1886 ( .A1(n2608), .A2(n2609), .ZN(n2607) );
OR_X1 U1887 ( .A1(n2528), .A2(n2610), .ZN(n2608) );
INV_X1 U1888 ( .A1(n2611), .ZN(n2606) );
INV_X1 U1889 ( .A1(n2577), .ZN(n2602) );
AND_X1 U1890 ( .A1(n2612), .A2(n2613), .ZN(n2537) );
NAND_X1 U1891 ( .A1(n2530), .A2(n2614), .ZN(n2613) );
NAND_X1 U1892 ( .A1(n2531), .A2(n2615), .ZN(n2614) );
INV_X1 U1893 ( .A1(n2532), .ZN(n2615) );
NOR_X1 U1894 ( .A1(n2471), .A2(n2616), .A3(n2527), .ZN(n2532) );
NAND_X1 U1895 ( .A1(n2362), .A2(n2617), .ZN(n2527) );
NAND_X1 U1896 ( .A1(n2618), .A2(n2528), .ZN(n2617) );
INV_X1 U1897 ( .A1(n2599), .ZN(n2618) );
AND_X1 U1898 ( .A1(n2412), .A2(n2528), .ZN(n2616) );
OR_X1 U1899 ( .A1(n2609), .A2(n2364), .ZN(n2531) );
NAND_X1 U1900 ( .A1(n2619), .A2(n2580), .ZN(n2612) );
INV_X1 U1901 ( .A1(n2605), .ZN(n2619) );
NOR_X1 U1902 ( .A1(n2620), .A2(n2621), .ZN(n2593) );
NOR_X1 U1903 ( .A1(n2520), .A2(n2622), .A3(n2521), .ZN(n2621) );
NOR_X1 U1904 ( .A1(n2471), .A2(n2508), .A3(n2412), .ZN(w1047) );
INV_X1 U1905 ( .A1(n2598), .ZN(n2520) );
NOR_X1 U1906 ( .A1(n2598), .A2(n2538), .ZN(n2620) );
NAND_X1 U1907 ( .A1(n2533), .A2(n2530), .ZN(n2538) );
INV_X1 U1908 ( .A1(n2508), .ZN(n2530) );
XOR_X1 U1909 ( .A1(n2611), .A2(n2623), .ZN(n2508) );
NOR_X1 U1910 ( .A1(n2624), .A2(n2580), .ZN(n2623) );
NOR_X1 U1911 ( .A1(n2471), .A2(n2412), .A3(n2521), .ZN(n2533) );
XOR_X1 U1912 ( .A1(n2625), .A2(n2626), .ZN(n2412) );
NOR_X1 U1913 ( .A1(n2627), .A2(n2362), .ZN(n2626) );
XOR_X1 U1914 ( .A1(n2610), .A2(n2628), .ZN(n2471) );
NOR_X1 U1915 ( .A1(n2629), .A2(n2362), .ZN(n2628) );
NOR_X1 U1916 ( .A1(n2625), .A2(n2611), .A3(n2577), .A4(n2610), .ZN(n2598) );
NAND_X1 U1917 ( .A1(n2609), .A2(n2630), .ZN(n2610) );
NAND_X1 U1918 ( .A1(n2631), .A2(n2632), .A3(n2629), .ZN(n2630) );
INV_X1 U1919 ( .A1(n2633), .ZN(n2629) );
NAND_X1 U1920 ( .A1(G200), .A2(n2634), .ZN(n2632) );
NAND_X1 U1921 ( .A1(n2635), .A2(G190), .ZN(n2631) );
NAND_X1 U1922 ( .A1(n2636), .A2(n2637), .A3(n2633), .ZN(n2609) );
NAND_X1 U1923 ( .A1(n2638), .A2(n2639), .A3(n2640), .A4(n2641), .ZN(n2633) );
OR_X1 U1924 ( .A1(n2642), .A2(n2448), .ZN(n2641) );
NAND_X1 U1925 ( .A1(n2643), .A2(n2448), .ZN(n2640) );
NAND_X1 U1926 ( .A1(n2644), .A2(G77), .ZN(n2639) );
NAND_X1 U1927 ( .A1(n2645), .A2(G50), .ZN(n2638) );
NAND_X1 U1928 ( .A1(n2635), .A2(n2646), .ZN(n2637) );
INV_X1 U1929 ( .A1(n2634), .ZN(n2635) );
NAND_X1 U1930 ( .A1(n2634), .A2(n2576), .ZN(n2636) );
NAND_X1 U1931 ( .A1(n2647), .A2(n2648), .A3(n2649), .ZN(n2634) );
NAND_X1 U1932 ( .A1(n2650), .A2(G238), .ZN(n2649) );
NAND_X1 U1933 ( .A1(n2651), .A2(n2652), .ZN(n2647) );
NAND_X1 U1934 ( .A1(n2653), .A2(n2654), .A3(n2655), .ZN(n2652) );
NAND_X1 U1935 ( .A1(G33), .A2(G97), .ZN(n2655) );
NAND_X1 U1936 ( .A1(n2656), .A2(G232), .ZN(n2654) );
NAND_X1 U1937 ( .A1(n2657), .A2(G226), .ZN(n2653) );
NAND_X1 U1938 ( .A1(n2601), .A2(n2658), .ZN(n2577) );
NAND_X1 U1939 ( .A1(n2659), .A2(n2660), .A3(n2579), .ZN(n2658) );
INV_X1 U1940 ( .A1(n2661), .ZN(n2579) );
NAND_X1 U1941 ( .A1(G200), .A2(n2662), .ZN(n2660) );
NAND_X1 U1942 ( .A1(n2663), .A2(G190), .ZN(n2659) );
NAND_X1 U1943 ( .A1(n2664), .A2(n2665), .A3(n2661), .ZN(n2601) );
NAND_X1 U1944 ( .A1(n2666), .A2(n2667), .A3(n2668), .A4(n2669), .ZN(n2661) );
NOR_X1 U1945 ( .A1(n2670), .A2(n2671), .ZN(n2669) );
NOR_X1 U1946 ( .A1(n2394), .A2(n2672), .ZN(n2671) );
INV_X1 U1947 ( .A1(G150), .ZN(n2394) );
NOR_X1 U1948 ( .A1(n2673), .A2(n2226), .ZN(n2670) );
NAND_X1 U1949 ( .A1(n2674), .A2(G68), .ZN(n2668) );
NAND_X1 U1950 ( .A1(n2675), .A2(n2228), .ZN(n2667) );
NAND_X1 U1951 ( .A1(G50), .A2(n2676), .ZN(n2666) );
NAND_X1 U1952 ( .A1(n2663), .A2(n2646), .ZN(n2665) );
INV_X1 U1953 ( .A1(n2662), .ZN(n2663) );
NAND_X1 U1954 ( .A1(n2662), .A2(n2576), .ZN(n2664) );
NAND_X1 U1955 ( .A1(n2677), .A2(n2648), .A3(n2678), .ZN(n2662) );
NAND_X1 U1956 ( .A1(n2650), .A2(G226), .ZN(n2678) );
NAND_X1 U1957 ( .A1(n2651), .A2(n2679), .ZN(n2677) );
NAND_X1 U1958 ( .A1(n2680), .A2(n2681), .A3(n2682), .ZN(n2679) );
NAND_X1 U1959 ( .A1(G33), .A2(G77), .ZN(n2682) );
NAND_X1 U1960 ( .A1(G223), .A2(n2656), .ZN(n2681) );
NAND_X1 U1961 ( .A1(G222), .A2(n2657), .ZN(n2680) );
NAND_X1 U1962 ( .A1(n2605), .A2(n2683), .ZN(n2611) );
NAND_X1 U1963 ( .A1(n2684), .A2(n2685), .A3(n2624), .ZN(n2683) );
INV_X1 U1964 ( .A1(n2686), .ZN(n2624) );
NAND_X1 U1965 ( .A1(G200), .A2(n2687), .ZN(n2685) );
NAND_X1 U1966 ( .A1(n2688), .A2(G190), .ZN(n2684) );
NAND_X1 U1967 ( .A1(n2689), .A2(n2690), .A3(n2686), .ZN(n2605) );
NAND_X1 U1968 ( .A1(n2691), .A2(n2692), .A3(n2693), .ZN(n2686) );
NOR_X1 U1969 ( .A1(n2694), .A2(n2695), .A3(n2696), .ZN(n2693) );
NOR_X1 U1970 ( .A1(n2226), .A2(n2642), .ZN(n2696) );
INV_X1 U1971 ( .A1(G58), .ZN(n2226) );
NOR_X1 U1972 ( .A1(G58), .A2(n2697), .ZN(n2695) );
NOR_X1 U1973 ( .A1(n2319), .A2(n2672), .ZN(n2694) );
INV_X1 U1974 ( .A1(G159), .ZN(n2319) );
NAND_X1 U1975 ( .A1(G68), .A2(n2698), .ZN(n2692) );
NAND_X1 U1976 ( .A1(n2699), .A2(n2700), .ZN(n2698) );
NAND_X1 U1977 ( .A1(n2674), .A2(G58), .ZN(n2700) );
NAND_X1 U1978 ( .A1(n2701), .A2(n2674), .ZN(n2691) );
NAND_X1 U1979 ( .A1(n2688), .A2(n2646), .ZN(n2690) );
INV_X1 U1980 ( .A1(n2687), .ZN(n2688) );
NAND_X1 U1981 ( .A1(n2687), .A2(n2576), .ZN(n2689) );
NAND_X1 U1982 ( .A1(n2702), .A2(n2648), .A3(n2703), .ZN(n2687) );
NAND_X1 U1983 ( .A1(n2650), .A2(G232), .ZN(n2703) );
NAND_X1 U1984 ( .A1(n2651), .A2(n2704), .ZN(n2702) );
NAND_X1 U1985 ( .A1(n2705), .A2(n2706), .A3(n2707), .ZN(n2704) );
NAND_X1 U1986 ( .A1(G33), .A2(G87), .ZN(n2707) );
NAND_X1 U1987 ( .A1(n2656), .A2(G226), .ZN(n2706) );
NAND_X1 U1988 ( .A1(G223), .A2(n2657), .ZN(n2705) );
NAND_X1 U1989 ( .A1(n2528), .A2(n2708), .ZN(n2625) );
NAND_X1 U1990 ( .A1(n2709), .A2(n2710), .A3(n2627), .ZN(n2708) );
INV_X1 U1991 ( .A1(n2711), .ZN(n2627) );
NAND_X1 U1992 ( .A1(G200), .A2(n2712), .ZN(n2710) );
NAND_X1 U1993 ( .A1(n2713), .A2(G190), .ZN(n2709) );
NAND_X1 U1994 ( .A1(n2714), .A2(n2715), .A3(n2711), .ZN(n2528) );
NAND_X1 U1995 ( .A1(n2716), .A2(n2717), .A3(n2718), .A4(n2719), .ZN(n2711) );
NAND_X1 U1996 ( .A1(n2675), .A2(n2440), .ZN(n2719) );
NAND_X1 U1997 ( .A1(G77), .A2(n2676), .ZN(n2718) );
NAND_X1 U1998 ( .A1(n2720), .A2(n2642), .ZN(n2676) );
NAND_X1 U1999 ( .A1(n2721), .A2(n2722), .ZN(n2642) );
NAND_X1 U2000 ( .A1(n2644), .A2(G87), .ZN(n2717) );
NAND_X1 U2001 ( .A1(n2645), .A2(G58), .ZN(n2716) );
NAND_X1 U2002 ( .A1(n2713), .A2(n2646), .ZN(n2715) );
INV_X1 U2003 ( .A1(n2712), .ZN(n2713) );
NAND_X1 U2004 ( .A1(n2712), .A2(n2576), .ZN(n2714) );
NAND_X1 U2005 ( .A1(n2723), .A2(n2648), .A3(n2724), .ZN(n2712) );
NAND_X1 U2006 ( .A1(n2650), .A2(G244), .ZN(n2724) );
NOR_X1 U2007 ( .A1(n2725), .A2(n2651), .ZN(n2650) );
NAND_X1 U2008 ( .A1(n2725), .A2(G274), .ZN(n2648) );
AND_X1 U2009 ( .A1(n2726), .A2(n2727), .ZN(n2725) );
NAND_X1 U2010 ( .A1(n2545), .A2(n2251), .ZN(n2727) );
NAND_X1 U2011 ( .A1(n2651), .A2(n2728), .ZN(n2723) );
NAND_X1 U2012 ( .A1(n2729), .A2(n2730), .A3(n2731), .ZN(n2728) );
NAND_X1 U2013 ( .A1(G107), .A2(G33), .ZN(n2731) );
NAND_X1 U2014 ( .A1(n2656), .A2(G238), .ZN(n2730) );
NAND_X1 U2015 ( .A1(n2657), .A2(G232), .ZN(n2729) );
NAND_X1 U2016 ( .A1(G116), .A2(n2732), .A3(n2733), .ZN(w1070) );
NAND_X1 U2017 ( .A1(n2734), .A2(n2735), .A3(n2736), .ZN(G364) );
NAND_X1 U2018 ( .A1(n2737), .A2(n2300), .ZN(n2736) );
OR_X1 U2019 ( .A1(n2265), .A2(n2300), .A3(n2726), .ZN(n2735) );
NOR_X1 U2020 ( .A1(n2738), .A2(G41), .ZN(n2300) );
NAND_X1 U2021 ( .A1(n2266), .A2(n2244), .A3(n2465), .A4(n2433), .ZN(n2265) );
NAND_X1 U2022 ( .A1(n2309), .A2(n2726), .ZN(n2734) );
NAND_X1 U2023 ( .A1(n2521), .A2(n2739), .ZN(n2309) );
NAND_X1 U2024 ( .A1(n2599), .A2(n2362), .ZN(n2739) );
NAND_X1 U2025 ( .A1(n2740), .A2(n2741), .ZN(n2599) );
NAND_X1 U2026 ( .A1(n2406), .A2(n2742), .ZN(n2741) );
NAND_X1 U2027 ( .A1(n2372), .A2(n2743), .ZN(n2742) );
NAND_X1 U2028 ( .A1(n2744), .A2(n2745), .ZN(n2743) );
NAND_X1 U2029 ( .A1(n2368), .A2(n2746), .ZN(n2745) );
OR_X1 U2030 ( .A1(n2363), .A2(n2365), .ZN(n2746) );
INV_X1 U2031 ( .A1(n2369), .ZN(n2744) );
INV_X1 U2032 ( .A1(n2747), .ZN(n2406) );
NAND_X1 U2033 ( .A1(n2748), .A2(n2749), .A3(G330), .ZN(n2521) );
NAND_X1 U2034 ( .A1(n2581), .A2(n2362), .ZN(n2749) );
INV_X1 U2035 ( .A1(n2364), .ZN(n2362) );
OR_X1 U2036 ( .A1(n2359), .A2(n2747), .A3(n2369), .A4(n2365), .ZN(n2581) );
NAND_X1 U2037 ( .A1(n2368), .A2(n2750), .ZN(n2365) );
NAND_X1 U2038 ( .A1(n2751), .A2(n2752), .A3(n2367), .ZN(n2750) );
INV_X1 U2039 ( .A1(n2753), .ZN(n2367) );
NAND_X1 U2040 ( .A1(G200), .A2(n2754), .ZN(n2752) );
NAND_X1 U2041 ( .A1(G190), .A2(n2755), .ZN(n2751) );
NAND_X1 U2042 ( .A1(n2756), .A2(n2757), .A3(n2753), .ZN(n2368) );
NAND_X1 U2043 ( .A1(n2758), .A2(n2759), .A3(n2760), .A4(n2761), .ZN(n2753) );
NAND_X1 U2044 ( .A1(n2762), .A2(G107), .ZN(n2761) );
NAND_X1 U2045 ( .A1(n2643), .A2(n2266), .ZN(n2760) );
NAND_X1 U2046 ( .A1(n2697), .A2(n2720), .ZN(n2643) );
NAND_X1 U2047 ( .A1(n2644), .A2(G116), .ZN(n2759) );
NAND_X1 U2048 ( .A1(n2645), .A2(G87), .ZN(n2758) );
NAND_X1 U2049 ( .A1(n2755), .A2(n2646), .ZN(n2757) );
NAND_X1 U2050 ( .A1(n2754), .A2(n2576), .ZN(n2756) );
NAND_X1 U2051 ( .A1(n2372), .A2(n2763), .ZN(n2369) );
NAND_X1 U2052 ( .A1(n2764), .A2(n2765), .A3(n2371), .ZN(n2763) );
INV_X1 U2053 ( .A1(n2766), .ZN(n2371) );
NAND_X1 U2054 ( .A1(G200), .A2(n2767), .ZN(n2765) );
NAND_X1 U2055 ( .A1(G190), .A2(n2768), .ZN(n2764) );
NAND_X1 U2056 ( .A1(n2769), .A2(n2770), .A3(n2766), .ZN(n2372) );
NAND_X1 U2057 ( .A1(n2771), .A2(n2772), .A3(n2773), .A4(n2774), .ZN(n2766) );
NOR_X1 U2058 ( .A1(n2775), .A2(n2776), .ZN(n2774) );
NOR_X1 U2059 ( .A1(n2440), .A2(n2672), .ZN(n2776) );
NOR_X1 U2060 ( .A1(n2699), .A2(n2266), .ZN(n2775) );
INV_X1 U2061 ( .A1(n2644), .ZN(n2699) );
OR_X1 U2062 ( .A1(n2732), .A2(n2720), .ZN(w1071) );
NAND_X1 U2063 ( .A1(n2675), .A2(n2433), .ZN(n2772) );
NAND_X1 U2064 ( .A1(n2762), .A2(G97), .ZN(n2771) );
INV_X1 U2065 ( .A1(n2777), .ZN(n2762) );
NAND_X1 U2066 ( .A1(n2768), .A2(n2646), .ZN(n2770) );
NAND_X1 U2067 ( .A1(n2767), .A2(n2576), .ZN(n2769) );
NAND_X1 U2068 ( .A1(n2740), .A2(n2778), .ZN(n2747) );
NAND_X1 U2069 ( .A1(n2779), .A2(n2780), .A3(n2408), .ZN(n2778) );
INV_X1 U2070 ( .A1(n2781), .ZN(n2408) );
NAND_X1 U2071 ( .A1(G200), .A2(n2782), .ZN(n2780) );
NAND_X1 U2072 ( .A1(G190), .A2(n2783), .ZN(n2779) );
NAND_X1 U2073 ( .A1(n2784), .A2(n2785), .A3(n2781), .ZN(n2740) );
NAND_X1 U2074 ( .A1(n2786), .A2(n2787), .A3(n2788), .A4(n2789), .ZN(n2781) );
NOR_X1 U2075 ( .A1(n2790), .A2(n2791), .ZN(n2789) );
NOR_X1 U2076 ( .A1(n2448), .A2(n2672), .ZN(n2791) );
INV_X1 U2077 ( .A1(n2645), .ZN(n2672) );
NOR_X1 U2078 ( .A1(n2673), .A2(n2433), .ZN(n2790) );
AND_X1 U2079 ( .A1(n2720), .A2(n2792), .ZN(n2673) );
OR_X1 U2080 ( .A1(n2721), .A2(n2389), .ZN(n2792) );
NAND_X1 U2081 ( .A1(n2674), .A2(G107), .ZN(n2788) );
NAND_X1 U2082 ( .A1(n2675), .A2(n2465), .ZN(n2787) );
INV_X1 U2083 ( .A1(G87), .ZN(n2465) );
NAND_X1 U2084 ( .A1(G87), .A2(n2793), .ZN(n2786) );
NAND_X1 U2085 ( .A1(n2783), .A2(n2646), .ZN(n2785) );
NAND_X1 U2086 ( .A1(n2782), .A2(n2576), .ZN(n2784) );
NAND_X1 U2087 ( .A1(n2363), .A2(n2794), .ZN(n2359) );
NAND_X1 U2088 ( .A1(n2795), .A2(n2796), .A3(n2361), .ZN(n2794) );
INV_X1 U2089 ( .A1(n2797), .ZN(n2361) );
NAND_X1 U2090 ( .A1(G200), .A2(n2798), .ZN(n2796) );
NAND_X1 U2091 ( .A1(G190), .A2(n2799), .ZN(n2795) );
NAND_X1 U2092 ( .A1(n2800), .A2(n2801), .A3(n2797), .ZN(n2363) );
NAND_X1 U2093 ( .A1(n2802), .A2(n2803), .A3(n2804), .A4(n2805), .ZN(n2797) );
NAND_X1 U2094 ( .A1(n2675), .A2(n2244), .ZN(n2805) );
NAND_X1 U2095 ( .A1(G116), .A2(n2793), .ZN(n2804) );
NAND_X1 U2096 ( .A1(n2777), .A2(n2720), .ZN(n2793) );
INV_X1 U2097 ( .A1(n2674), .ZN(n2720) );
NOR_X1 U2098 ( .A1(n2721), .A2(n2543), .ZN(n2674) );
NAND_X1 U2099 ( .A1(n2721), .A2(n2697), .A3(n2806), .ZN(n2777) );
NAND_X1 U2100 ( .A1(G33), .A2(n2726), .ZN(n2806) );
INV_X1 U2101 ( .A1(n2675), .ZN(n2697) );
NOR_X1 U2102 ( .A1(n2722), .A2(n2586), .ZN(n2675) );
NAND_X1 U2103 ( .A1(G20), .A2(n2726), .ZN(n2722) );
NAND_X1 U2104 ( .A1(n2644), .A2(G283), .ZN(n2803) );
NOR_X1 U2105 ( .A1(n2389), .A2(G20), .A3(n2721), .ZN(n2644) );
NAND_X1 U2106 ( .A1(n2645), .A2(G97), .ZN(n2802) );
NOR_X1 U2107 ( .A1(G20), .A2(G33), .A3(n2721), .ZN(n2645) );
NAND_X1 U2108 ( .A1(n2807), .A2(n2405), .A3(G1), .ZN(n2721) );
NAND_X1 U2109 ( .A1(n2389), .A2(n2586), .ZN(n2405) );
INV_X1 U2110 ( .A1(G33), .ZN(n2389) );
NAND_X1 U2111 ( .A1(n2586), .A2(n2543), .ZN(n2807) );
NAND_X1 U2112 ( .A1(n2799), .A2(n2646), .ZN(n2801) );
NAND_X1 U2113 ( .A1(n2798), .A2(n2576), .ZN(n2800) );
INV_X1 U2114 ( .A1(G169), .ZN(n2576) );
NAND_X1 U2115 ( .A1(n2808), .A2(n2364), .ZN(n2748) );
NOR_X1 U2116 ( .A1(n2185), .A2(n2580), .ZN(n2364) );
NAND_X1 U2117 ( .A1(G213), .A2(G13), .A3(n2726), .A4(n2543), .ZN(n2580) );
INV_X1 U2118 ( .A1(G20), .ZN(n2543) );
INV_X1 U2119 ( .A1(G1), .ZN(n2726) );
INV_X1 U2120 ( .A1(G343), .ZN(n2185) );
NAND_X1 U2121 ( .A1(n2809), .A2(n2810), .ZN(n2808) );
NAND_X1 U2122 ( .A1(G179), .A2(n2811), .ZN(n2810) );
NAND_X1 U2123 ( .A1(n2799), .A2(n2768), .A3(n2783), .A4(n2755), .ZN(n2811) );
INV_X1 U2124 ( .A1(n2754), .ZN(n2755) );
INV_X1 U2125 ( .A1(n2782), .ZN(n2783) );
INV_X1 U2126 ( .A1(n2767), .ZN(n2768) );
INV_X1 U2127 ( .A1(n2798), .ZN(n2799) );
NAND_X1 U2128 ( .A1(n2812), .A2(n2646), .ZN(n2809) );
INV_X1 U2129 ( .A1(G179), .ZN(n2646) );
NAND_X1 U2130 ( .A1(n2754), .A2(n2767), .A3(n2782), .A4(n2798), .ZN(n2812) );
NAND_X1 U2131 ( .A1(n2813), .A2(n2814), .A3(n2815), .ZN(n2798) );
NAND_X1 U2132 ( .A1(n2651), .A2(n2816), .ZN(n2815) );
NAND_X1 U2133 ( .A1(n2817), .A2(n2818), .A3(n2819), .ZN(n2816) );
NAND_X1 U2134 ( .A1(G303), .A2(G33), .ZN(n2819) );
NAND_X1 U2135 ( .A1(n2656), .A2(G264), .ZN(n2818) );
NAND_X1 U2136 ( .A1(n2657), .A2(G257), .ZN(n2817) );
NAND_X1 U2137 ( .A1(G270), .A2(n2820), .ZN(n2813) );
NAND_X1 U2138 ( .A1(n2821), .A2(n2822), .A3(n2823), .ZN(n2782) );
NAND_X1 U2139 ( .A1(G274), .A2(n2824), .ZN(n2823) );
OR_X1 U2140 ( .A1(n2825), .A2(n2824), .A3(n2651), .ZN(n2822) );
NAND_X1 U2141 ( .A1(n2651), .A2(n2826), .ZN(n2821) );
NAND_X1 U2142 ( .A1(n2827), .A2(n2828), .A3(n2829), .ZN(n2826) );
NAND_X1 U2143 ( .A1(G116), .A2(G33), .ZN(n2829) );
NAND_X1 U2144 ( .A1(n2656), .A2(G244), .ZN(n2828) );
NAND_X1 U2145 ( .A1(n2657), .A2(G238), .ZN(n2827) );
NAND_X1 U2146 ( .A1(n2830), .A2(n2814), .A3(n2831), .ZN(n2767) );
NAND_X1 U2147 ( .A1(n2651), .A2(n2832), .ZN(n2831) );
NAND_X1 U2148 ( .A1(n2833), .A2(n2834), .A3(n2835), .ZN(n2832) );
NAND_X1 U2149 ( .A1(G283), .A2(G33), .ZN(n2835) );
NAND_X1 U2150 ( .A1(G250), .A2(n2656), .ZN(n2834) );
NAND_X1 U2151 ( .A1(n2657), .A2(G244), .ZN(n2833) );
NAND_X1 U2152 ( .A1(G257), .A2(n2820), .ZN(n2830) );
NAND_X1 U2153 ( .A1(n2836), .A2(n2814), .A3(n2837), .ZN(n2754) );
NAND_X1 U2154 ( .A1(n2651), .A2(n2838), .ZN(n2837) );
NAND_X1 U2155 ( .A1(n2839), .A2(n2840), .A3(n2841), .ZN(n2838) );
NAND_X1 U2156 ( .A1(G294), .A2(G33), .ZN(n2841) );
NAND_X1 U2157 ( .A1(G257), .A2(n2656), .ZN(n2840) );
NOR_X1 U2158 ( .A1(n2657), .A2(G33), .ZN(n2656) );
NAND_X1 U2159 ( .A1(G250), .A2(n2657), .ZN(n2839) );
NOR_X1 U2160 ( .A1(G33), .A2(G1698), .ZN(n2657) );
NAND_X1 U2161 ( .A1(G274), .A2(n2842), .ZN(n2814) );
NAND_X1 U2162 ( .A1(G264), .A2(n2820), .ZN(n2836) );
NOR_X1 U2163 ( .A1(n2842), .A2(n2651), .ZN(n2820) );
AND_X1 U2164 ( .A1(G1), .A2(n2843), .A3(G13), .ZN(n2651) );
NAND_X1 U2165 ( .A1(G41), .A2(G33), .ZN(n2843) );
AND_X1 U2166 ( .A1(n2824), .A2(n2545), .ZN(n2842) );
INV_X1 U2167 ( .A1(G41), .ZN(n2545) );
NOR_X1 U2168 ( .A1(n2251), .A2(G1), .ZN(n2824) );
INV_X1 U2169 ( .A1(G45), .ZN(n2251) );
NOR_X1 U2170 ( .A1(n2844), .A2(n2845), .A3(n2846), .ZN(G361) );
NOR_X1 U2171 ( .A1(n2738), .A2(n2847), .A3(n2825), .ZN(n2846) );
INV_X1 U2172 ( .A1(G250), .ZN(n2825) );
NOR_X1 U2173 ( .A1(G257), .A2(G264), .ZN(n2847) );
NOR_X1 U2174 ( .A1(n2388), .A2(n2733), .A3(n2848), .ZN(n2845) );
NOR_X1 U2175 ( .A1(n2849), .A2(n2850), .ZN(n2848) );
NAND_X1 U2176 ( .A1(n2851), .A2(n2852), .A3(n2853), .A4(n2854), .ZN(n2850) );
NAND_X1 U2177 ( .A1(G238), .A2(G68), .ZN(n2854) );
NAND_X1 U2178 ( .A1(G244), .A2(G77), .ZN(n2853) );
NAND_X1 U2179 ( .A1(G250), .A2(G87), .ZN(n2852) );
NAND_X1 U2180 ( .A1(G257), .A2(G97), .ZN(n2851) );
NAND_X1 U2181 ( .A1(n2855), .A2(n2856), .A3(n2857), .A4(n2858), .ZN(n2849) );
NAND_X1 U2182 ( .A1(G264), .A2(G107), .ZN(n2858) );
NAND_X1 U2183 ( .A1(G270), .A2(G116), .ZN(n2857) );
NAND_X1 U2184 ( .A1(G226), .A2(G50), .ZN(n2856) );
NAND_X1 U2185 ( .A1(G232), .A2(G58), .ZN(n2855) );
INV_X1 U2186 ( .A1(n2592), .ZN(n2733) );
INV_X1 U2187 ( .A1(n2738), .ZN(n2388) );
NAND_X1 U2188 ( .A1(G1), .A2(n2586), .A3(G20), .ZN(n2738) );
INV_X1 U2189 ( .A1(G13), .ZN(n2586) );
NOR_X1 U2190 ( .A1(n2252), .A2(n2592), .ZN(n2844) );
NAND_X1 U2191 ( .A1(G20), .A2(G1), .A3(G13), .ZN(n2592) );
INV_X1 U2192 ( .A1(n2737), .ZN(n2252) );
NOR_X1 U2193 ( .A1(n2228), .A2(n2701), .ZN(n2737) );
XOR_X1 U2194 ( .A1(n2404), .A2(n2272), .ZN(w1061) );
XNOR_X1 U2195 ( .A1(n2859), .A2(n2860), .ZN(w1052) );
XOR_X1 U2196 ( .A1(w1056), .A2(w1057), .ZN(n2860) );
XNOR_X1 U2197 ( .A1(w1058), .A2(w1059), .ZN(n2859) );
XOR_X1 U2198 ( .A1(n2861), .A2(n2862), .ZN(w1053) );
XOR_X1 U2199 ( .A1(w1062), .A2(w1063), .ZN(n2862) );
XNOR_X1 U2200 ( .A1(w1064), .A2(w1065), .ZN(n2861) );
NAND_X1 U2201 ( .A1(G87), .A2(n2863), .ZN(G355) );
NAND_X1 U2202 ( .A1(n2266), .A2(n2433), .ZN(n2863) );
AND_X1 U2203 ( .A1(n2701), .A2(n2440), .A3(n2228), .ZN(G353) );
NOR_X1 U2204 ( .A1(G58), .A2(G68), .ZN(n2701) );
XOR_X1 U2205 ( .A1(n2250), .A2(n2337), .ZN(w1069) );
XNOR_X1 U2206 ( .A1(n2864), .A2(n2732), .ZN(w1073) );
XOR_X1 U2207 ( .A1(n2266), .A2(n2433), .ZN(n2732) );
INV_X1 U2208 ( .A1(G97), .ZN(n2433) );
INV_X1 U2209 ( .A1(G107), .ZN(n2266) );
XOR_X1 U2210 ( .A1(n2244), .A2(w1072), .ZN(n2864) );
INV_X1 U2211 ( .A1(G116), .ZN(n2244) );
NAND_X1 U2212 ( .A1(n2865), .A2(n2866), .A3(n2867), .ZN(w1067) );
NAND_X1 U2213 ( .A1(n2271), .A2(n2868), .ZN(n2867) );
INV_X1 U2214 ( .A1(n2869), .ZN(w1077) );
NOR_X1 U2215 ( .A1(n2440), .A2(n2448), .ZN(n2271) );
NAND_X1 U2216 ( .A1(n2869), .A2(n2448), .A3(G77), .ZN(n2866) );
NAND_X1 U2217 ( .A1(n2870), .A2(n2440), .ZN(w1074) );
INV_X1 U2218 ( .A1(G77), .ZN(n2440) );
XOR_X1 U2219 ( .A1(n2448), .A2(n2869), .ZN(n2870) );
XNOR_X1 U2220 ( .A1(n2228), .A2(w1076), .ZN(w1075) );
INV_X1 U2221 ( .A1(G50), .ZN(n2228) );
INV_X1 U2222 ( .A1(G68), .ZN(n2448) );
XOR_X1 X1000 ( .A1(w1000), .A2(KEYINPUT0), .ZN(n2178) );
XNOR_X1 X1001 ( .A1(w1001), .A2(KEYINPUT1), .ZN(n2177) );
XOR_X1 X1002 ( .A1(w1002), .A2(KEYINPUT2), .ZN(G405) );
XNOR_X1 X1003 ( .A1(w1003), .A2(KEYINPUT3), .ZN(n2180) );
XOR_X1 X1004 ( .A1(w1004), .A2(KEYINPUT4), .ZN(n2186) );
XNOR_X1 X1005 ( .A1(w1005), .A2(KEYINPUT5), .ZN(G375) );
XOR_X1 X1006 ( .A1(w1006), .A2(KEYINPUT6), .ZN(G402) );
XNOR_X1 X1007 ( .A1(w1007), .A2(KEYINPUT7), .ZN(n2173) );
XOR_X1 X1008 ( .A1(w1008), .A2(KEYINPUT8), .ZN(w1000) );
XNOR_X1 X1009 ( .A1(w1009), .A2(KEYINPUT9), .ZN(w1004) );
XOR_X1 X1010 ( .A1(w1010), .A2(KEYINPUT10), .ZN(n2179) );
XNOR_X1 X1011 ( .A1(w1011), .A2(KEYINPUT11), .ZN(n2189) );
XOR_X1 X1012 ( .A1(w1012), .A2(KEYINPUT12), .ZN(n2188) );
XNOR_X1 X1013 ( .A1(w1013), .A2(KEYINPUT13), .ZN(G387) );
XOR_X1 X1014 ( .A1(w1014), .A2(KEYINPUT14), .ZN(w1010) );
XNOR_X1 X1015 ( .A1(w1015), .A2(KEYINPUT15), .ZN(n2190) );
XOR_X1 X1016 ( .A1(w1016), .A2(KEYINPUT16), .ZN(n2187) );
XNOR_X1 X1017 ( .A1(w1017), .A2(KEYINPUT17), .ZN(G393) );
XOR_X1 X1018 ( .A1(G330), .A2(KEYINPUT18), .ZN(w1018) );
XNOR_X1 X1019 ( .A1(w1019), .A2(KEYINPUT19), .ZN(n2192) );
XOR_X1 X1020 ( .A1(w1020), .A2(KEYINPUT20), .ZN(n2256) );
XNOR_X1 X1021 ( .A1(w1021), .A2(KEYINPUT21), .ZN(n2340) );
XOR_X1 X1022 ( .A1(w1022), .A2(KEYINPUT22), .ZN(n2305) );
XNOR_X1 X1023 ( .A1(w1023), .A2(KEYINPUT23), .ZN(n2342) );
XOR_X1 X1024 ( .A1(w1024), .A2(KEYINPUT24), .ZN(n2344) );
XNOR_X1 X1025 ( .A1(w1025), .A2(KEYINPUT25), .ZN(n2351) );
XOR_X1 X1026 ( .A1(w1026), .A2(KEYINPUT26), .ZN(n2196) );
XNOR_X1 X1027 ( .A1(w1027), .A2(KEYINPUT27), .ZN(n2195) );
XOR_X1 X1028 ( .A1(w1028), .A2(KEYINPUT28), .ZN(n2258) );
XNOR_X1 X1029 ( .A1(w1029), .A2(KEYINPUT29), .ZN(n2349) );
XOR_X1 X1030 ( .A1(w1030), .A2(KEYINPUT30), .ZN(n2310) );
XNOR_X1 X1031 ( .A1(w1031), .A2(KEYINPUT31), .ZN(n2350) );
XOR_X1 X1032 ( .A1(w1032), .A2(KEYINPUT32), .ZN(n2345) );
XNOR_X1 X1033 ( .A1(w1033), .A2(KEYINPUT33), .ZN(n2373) );
XOR_X1 X1034 ( .A1(w1034), .A2(KEYINPUT34), .ZN(n2410) );
XNOR_X1 X1035 ( .A1(w1035), .A2(KEYINPUT35), .ZN(n2301) );
XOR_X1 X1036 ( .A1(w1036), .A2(KEYINPUT36), .ZN(n2478) );
XNOR_X1 X1037 ( .A1(w1037), .A2(KEYINPUT37), .ZN(n2512) );
XOR_X1 X1038 ( .A1(w1038), .A2(KEYINPUT38), .ZN(n2514) );
XNOR_X1 X1039 ( .A1(w1039), .A2(KEYINPUT39), .ZN(n2535) );
XOR_X1 X1040 ( .A1(w1040), .A2(KEYINPUT40), .ZN(n2515) );
XNOR_X1 X1041 ( .A1(w1041), .A2(KEYINPUT41), .ZN(n2539) );
XOR_X1 X1042 ( .A1(w1042), .A2(KEYINPUT42), .ZN(n2583) );
XNOR_X1 X1043 ( .A1(w1043), .A2(KEYINPUT43), .ZN(n2594) );
XOR_X1 X1044 ( .A1(w1044), .A2(KEYINPUT44), .ZN(n2590) );
XNOR_X1 X1045 ( .A1(w1045), .A2(KEYINPUT45), .ZN(n2518) );
XOR_X1 X1046 ( .A1(w1046), .A2(KEYINPUT46), .ZN(n2482) );
XNOR_X1 X1047 ( .A1(w1047), .A2(KEYINPUT47), .ZN(n2622) );
XOR_X1 X1048 ( .A1(w1048), .A2(KEYINPUT48), .ZN(n2411) );
XNOR_X1 X1049 ( .A1(w1049), .A2(KEYINPUT49), .ZN(n2413) );
XOR_X1 X1050 ( .A1(w1050), .A2(KEYINPUT50), .ZN(n2445) );
XNOR_X1 X1051 ( .A1(w1051), .A2(KEYINPUT51), .ZN(n2523) );
XOR_X1 X1052 ( .A1(w1052), .A2(KEYINPUT52), .ZN(n2272) );
XNOR_X1 X1053 ( .A1(w1053), .A2(KEYINPUT53), .ZN(n2404) );
XOR_X1 X1054 ( .A1(w1054), .A2(KEYINPUT54), .ZN(n2268) );
XNOR_X1 X1055 ( .A1(w1055), .A2(KEYINPUT55), .ZN(G358) );
XOR_X1 X1056 ( .A1(G244), .A2(KEYINPUT56), .ZN(w1056) );
XNOR_X1 X1057 ( .A1(G238), .A2(KEYINPUT57), .ZN(w1057) );
XOR_X1 X1058 ( .A1(G226), .A2(KEYINPUT58), .ZN(w1058) );
XNOR_X1 X1059 ( .A1(G232), .A2(KEYINPUT59), .ZN(w1059) );
XOR_X1 X1060 ( .A1(w1060), .A2(KEYINPUT60), .ZN(n2401) );
XNOR_X1 X1061 ( .A1(w1061), .A2(KEYINPUT61), .ZN(w1055) );
XOR_X1 X1062 ( .A1(G257), .A2(KEYINPUT62), .ZN(w1062) );
XNOR_X1 X1063 ( .A1(G250), .A2(KEYINPUT63), .ZN(w1063) );
XOR_X1 X1064 ( .A1(G270), .A2(KEYINPUT64), .ZN(w1064) );
XNOR_X1 X1065 ( .A1(G264), .A2(KEYINPUT65), .ZN(w1065) );
XOR_X1 X1066 ( .A1(w1066), .A2(KEYINPUT66), .ZN(n2337) );
XNOR_X1 X1067 ( .A1(w1067), .A2(KEYINPUT67), .ZN(n2250) );
XOR_X1 X1068 ( .A1(w1068), .A2(KEYINPUT68), .ZN(n2335) );
XNOR_X1 X1069 ( .A1(w1069), .A2(KEYINPUT69), .ZN(G351) );
XOR_X1 X1070 ( .A1(w1070), .A2(KEYINPUT70), .ZN(n2582) );
XNOR_X1 X1071 ( .A1(w1071), .A2(KEYINPUT71), .ZN(n2773) );
XOR_X1 X1072 ( .A1(G87), .A2(KEYINPUT72), .ZN(w1072) );
XNOR_X1 X1073 ( .A1(w1073), .A2(KEYINPUT73), .ZN(w1066) );
XOR_X1 X1074 ( .A1(w1074), .A2(KEYINPUT74), .ZN(n2865) );
XNOR_X1 X1075 ( .A1(w1075), .A2(KEYINPUT75), .ZN(n2869) );
XOR_X1 X1076 ( .A1(G58), .A2(KEYINPUT76), .ZN(w1076) );
XNOR_X1 X1077 ( .A1(w1077), .A2(KEYINPUT77), .ZN(n2868) );
