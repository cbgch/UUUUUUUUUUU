module s208(
    P_0,
    C_8,
    C_7,
    C_6,
    C_5,
    C_4,
    C_3,
    C_2,
    C_1,
    C_0,
    Z);
    input P_0;
    input C_8;
    input C_7;
    input C_6;
    input C_5;
    input C_4;
    input C_3;
    input C_2;
    input C_1;
    input C_0;
    output Z;

    // Internal wires
    wire X_4;
    wire X_3;
    wire X_2;
    wire X_1;
    wire X_8;
    wire X_7;
    wire X_6;
    wire X_5;
    wire I73_1;
    wire I73_2;
    wire I7_1;
    wire I7_2;
    wire I88_1;
    wire I88_2;
    wire I48;
    wire I49;
    wire I50;
    wire I68;
    wire I105_1;
    wire I105_2;
    wire I182_1;
    wire I182_2;
    wire I148;
    wire I149;
    wire I161;
    wire I164;
    wire I212;
    wire I213;
    wire I214;
    wire I215;
    wire I216;
    wire I225;
    wire I240;
    wire I241;
    wire I242;
    wire I243;
    wire I244;
    wire I252;
    wire I282;
    wire I283;
    wire I286;
    wire I287;
    wire I306;
    wire I307;
    wire I310;
    wire I311;
    wire I73_3;
    wire I73_4;
    wire I7_3;
    wire I7_4;
    wire I88_3;
    wire I88_4;
    wire I105_3;
    wire I105_4;
    wire I182_3;
    wire I182_4;
    wire I191_1;
    wire I1_2;
    wire P_5;
    wire P_6;
    wire P_7;
    wire P_8;
    wire I295_1;
    wire I295_2;
    wire I319_1;
    wire I319_2;
    wire I270_3;
    wire I70_1;
    wire I13;
    wire I15;
    wire I95_1;
    wire I167_1;
    wire I170_1;
    wire I113;
    wire I188_1;
    wire I291_1;
    wire I291_2;
    wire I315_1;
    wire I315_2;
    wire I270_2;
    wire I12;
    wire I62;
    wire I64;
    wire I66;
    wire I110;
    wire I111;
    wire I159;
    wire I163;
    wire I165;
    wire I222;
    wire I224;
    wire I249;
    wire I251;
    wire I269_1;
    wire I269_2;
    wire I14;
    wire I2_1;
    wire I69;
    wire I112;
    wire I162;
    wire P_1;
    wire P_2;
    wire P_3;
    wire P_4;
    wire I209_1;
    wire I205_2;
    wire I206_2;
    wire I207_2;
    wire I208_2;
    wire I290;
    wire I314;
    DFFSRX1 g_X_4 (.D(I12),.Q(X_4),.CK(clk), .SN(setn), .RN(1'b1), .QN());
    DFFSRX1 g_X_3 (.D(I13),.Q(X_3),.CK(clk), .SN(setn), .RN(1'b1), .QN());
    DFFSRX1 g_X_2 (.D(I14),.Q(X_2),.CK(clk), .SN(setn), .RN(1'b1), .QN());
    DFFSRX1 g_X_1 (.D(I15),.Q(X_1),.CK(clk), .SN(setn), .RN(1'b1), .QN());
    DFFSRX1 g_X_8 (.D(I110),.Q(X_8),.CK(clk), .RN(rstn), .SN(1'b1), .QN());
    DFFSRX1 g_X_7 (.D(I111),.Q(X_7),.CK(clk), .RN(rstn), .SN(1'b1), .QN());
    DFFSRX1 g_X_6 (.D(I112),.Q(X_6),.CK(clk), .SN(setn), .RN(1'b1), .QN());
    DFFSRX1 g_X_5 (.D(I113),.Q(X_5),.CK(clk), .SN(setn), .RN(1'b1), .QN());
    INVX1 g_I73_1 (.A(I69),.Y(I73_1));
    INVX1 g_I73_2 (.A(X_3),.Y(I73_2));
    INVX1 g_I7_1 (.A(I66),.Y(I7_1));
    INVX1 g_I7_2 (.A(X_2),.Y(I7_2));
    INVX1 g_I88_1 (.A(X_1),.Y(I88_1));
    INVX1 g_I88_2 (.A(P_0),.Y(I88_2));
    INVX1 g_I48 (.A(P_0),.Y(I48));
    INVX1 g_I49 (.A(X_4),.Y(I49));
    INVX1 g_I50 (.A(X_3),.Y(I50));
    INVX1 g_I68 (.A(I69),.Y(I68));
    INVX1 g_I105_1 (.A(I163),.Y(I105_1));
    INVX1 g_I105_2 (.A(X_6),.Y(I105_2));
    INVX1 g_I182_1 (.A(X_5),.Y(I182_1));
    INVX1 g_I182_2 (.A(I1_2),.Y(I182_2));
    INVX1 g_I148 (.A(X_7),.Y(I148));
    INVX1 g_I149 (.A(X_6),.Y(I149));
    INVX1 g_I161 (.A(I162),.Y(I161));
    INVX1 g_I164 (.A(I163),.Y(I164));
    INVX1 g_I212 (.A(P_0),.Y(I212));
    INVX1 g_I213 (.A(X_1),.Y(I213));
    INVX1 g_I214 (.A(X_2),.Y(I214));
    INVX1 g_I215 (.A(X_3),.Y(I215));
    INVX1 g_I216 (.A(X_4),.Y(I216));
    INVX1 g_I225 (.A(I224),.Y(I225));
    INVX1 g_I240 (.A(P_0),.Y(I240));
    INVX1 g_I241 (.A(X_5),.Y(I241));
    INVX1 g_I242 (.A(X_6),.Y(I242));
    INVX1 g_I243 (.A(X_7),.Y(I243));
    INVX1 g_I244 (.A(X_8),.Y(I244));
    INVX1 g_I252 (.A(I251),.Y(I252));
    INVX1 g_I282 (.A(P_2),.Y(I282));
    INVX1 g_I283 (.A(P_3),.Y(I283));
    INVX1 g_I286 (.A(C_2),.Y(I286));
    INVX1 g_I287 (.A(C_3),.Y(I287));
    INVX1 g_I306 (.A(P_6),.Y(I306));
    INVX1 g_I307 (.A(P_7),.Y(I307));
    INVX1 g_I310 (.A(C_6),.Y(I310));
    INVX1 g_I311 (.A(C_7),.Y(I311));
    AND2X1 g_I73_3 (.A(I69),.B(I73_2),.Y(I73_3));
    AND2X1 g_I73_4 (.A(X_3),.B(I73_1),.Y(I73_4));
    AND2X1 g_I7_3 (.A(I66),.B(I7_2),.Y(I7_3));
    AND2X1 g_I7_4 (.A(X_2),.B(I7_1),.Y(I7_4));
    AND2X1 g_I88_3 (.A(X_1),.B(I88_2),.Y(I88_3));
    AND2X1 g_I88_4 (.A(P_0),.B(I88_1),.Y(I88_4));
    AND2X1 g_I105_3 (.A(I163),.B(I105_2),.Y(I105_3));
    AND2X1 g_I105_4 (.A(X_6),.B(I105_1),.Y(I105_4));
    AND2X1 g_I182_3 (.A(X_5),.B(I182_2),.Y(I182_3));
    AND2X1 g_I182_4 (.A(I1_2),.B(I182_1),.Y(I182_4));
    AND2X1 g_I191_1 (.A(I164),.B(X_6),.Y(I191_1));
    AND2X1 g_I1_2 (.A(I2_1),.B(P_0),.Y(I1_2));
    AND2X1 g_P_5 (.A(I209_1),.B(I205_2),.Y(P_5));
    AND2X1 g_P_6 (.A(I209_1),.B(I206_2),.Y(P_6));
    AND2X1 g_P_7 (.A(I209_1),.B(I207_2),.Y(P_7));
    AND2X1 g_P_8 (.A(I209_1),.B(I208_2),.Y(P_8));
    AND2X1 g_I295_1 (.A(P_1),.B(C_1),.Y(I295_1));
    AND2X1 g_I295_2 (.A(P_0),.B(C_0),.Y(I295_2));
    AND2X1 g_I319_1 (.A(P_5),.B(C_5),.Y(I319_1));
    AND2X1 g_I319_2 (.A(P_4),.B(C_4),.Y(I319_2));
    AND2X1 g_I270_3 (.A(P_8),.B(C_8),.Y(I270_3));
    OR3X1 g_I70_1 (.A(I68),.B(X_4),.C(I50),.Y(I70_1));
    OR2X1 g_I13 (.A(I73_3),.B(I73_4),.Y(I13));
    OR2X1 g_I15 (.A(I88_3),.B(I88_4),.Y(I15));
    OR3X1 g_I95_1 (.A(I64),.B(I50),.C(I48),.Y(I95_1));
    OR3X1 g_I167_1 (.A(I165),.B(X_8),.C(I148),.Y(I167_1));
    OR2X1 g_I170_1 (.A(I165),.B(X_7),.Y(I170_1));
    OR2X1 g_I113 (.A(I182_3),.B(I182_4),.Y(I113));
    OR3X1 g_I188_1 (.A(I163),.B(I149),.C(I148),.Y(I188_1));
    OR2X1 g_I291_1 (.A(I283),.B(I287),.Y(I291_1));
    OR2X1 g_I291_2 (.A(I282),.B(I286),.Y(I291_2));
    OR2X1 g_I315_1 (.A(I307),.B(I311),.Y(I315_1));
    OR2X1 g_I315_2 (.A(I306),.B(I310),.Y(I315_2));
    OR2X1 g_I270_2 (.A(I269_1),.B(I269_2),.Y(I270_2));
    OR2X1 g_Z (.A(I270_2),.B(I270_3),.Y(Z));
    NAND2X1 g_I12 (.A(I70_1),.B(I62),.Y(I12));
    NAND2X1 g_I62 (.A(I95_1),.B(X_4),.Y(I62));
    NAND2X1 g_I64 (.A(X_1),.B(X_2),.Y(I64));
    NAND2X1 g_I66 (.A(X_1),.B(P_0),.Y(I66));
    NAND2X1 g_I110 (.A(I167_1),.B(I159),.Y(I110));
    NAND2X1 g_I111 (.A(I170_1),.B(I161),.Y(I111));
    NAND2X1 g_I159 (.A(I188_1),.B(X_8),.Y(I159));
    NAND2X1 g_I163 (.A(X_5),.B(I1_2),.Y(I163));
    NAND2X1 g_I165 (.A(I164),.B(X_6),.Y(I165));
    NAND2X1 g_I222 (.A(I225),.B(I214),.Y(I222));
    NAND2X1 g_I224 (.A(I213),.B(P_0),.Y(I224));
    NAND2X1 g_I249 (.A(I252),.B(I242),.Y(I249));
    NAND2X1 g_I251 (.A(I241),.B(P_0),.Y(I251));
    NAND3X1 g_I269_1 (.A(I291_1),.B(I291_2),.C(I290),.Y(I269_1));
    NAND3X1 g_I269_2 (.A(I315_1),.B(I315_2),.C(I314),.Y(I269_2));
    NOR2X1 g_I14 (.A(I7_3),.B(I7_4),.Y(I14));
    NOR3X1 g_I2_1 (.A(I64),.B(I49),.C(I50),.Y(I2_1));
    NOR2X1 g_I69 (.A(I64),.B(I48),.Y(I69));
    NOR2X1 g_I112 (.A(I105_3),.B(I105_4),.Y(I112));
    NOR2X1 g_I162 (.A(I148),.B(I191_1),.Y(I162));
    NOR2X1 g_P_1 (.A(I212),.B(I213),.Y(P_1));
    NOR2X1 g_P_2 (.A(I214),.B(I224),.Y(P_2));
    NOR2X1 g_P_3 (.A(I215),.B(I222),.Y(P_3));
    NOR3X1 g_P_4 (.A(X_3),.B(I222),.C(I216),.Y(P_4));
    NOR4X1 g_I209_1 (.A(X_4),.B(X_2),.C(X_3),.D(X_1),.Y(I209_1));
    NOR2X1 g_I205_2 (.A(I240),.B(I241),.Y(I205_2));
    NOR2X1 g_I206_2 (.A(I242),.B(I251),.Y(I206_2));
    NOR2X1 g_I207_2 (.A(I243),.B(I249),.Y(I207_2));
    NOR3X1 g_I208_2 (.A(X_7),.B(I249),.C(I244),.Y(I208_2));
    NOR2X1 g_I290 (.A(I295_1),.B(I295_2),.Y(I290));
    NOR2X1 g_I314 (.A(I319_1),.B(I319_2),.Y(I314));
    
endmodule