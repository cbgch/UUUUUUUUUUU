module c1908 ( G953,G898,G224,G902,G952,G214,G900,G221,G110,G217,G119,G137,G128,G234,
G472,G101,G210,G237,G125,G122,G113,G116,G469,G140,G227,G107,G104,G134,
G131,G146,G475,G143,G478,KEYINPUT0,KEYINPUT1,KEYINPUT2,KEYINPUT3,KEYINPUT4,KEYINPUT5,KEYINPUT6,KEYINPUT7,KEYINPUT8,
KEYINPUT9,KEYINPUT10,KEYINPUT11,KEYINPUT12,KEYINPUT13,KEYINPUT14,KEYINPUT15,KEYINPUT16,KEYINPUT17,KEYINPUT18,KEYINPUT19,KEYINPUT20,KEYINPUT21,KEYINPUT22,
KEYINPUT23,KEYINPUT24,KEYINPUT25,KEYINPUT26,KEYINPUT27,KEYINPUT28,KEYINPUT29,KEYINPUT30,KEYINPUT31,KEYINPUT32,KEYINPUT33,KEYINPUT34,KEYINPUT35,KEYINPUT36,
KEYINPUT37,KEYINPUT38,KEYINPUT39,KEYINPUT40,KEYINPUT41,KEYINPUT42,KEYINPUT43,KEYINPUT44,KEYINPUT45,KEYINPUT46,KEYINPUT47,KEYINPUT48,KEYINPUT49,KEYINPUT50,
KEYINPUT51,KEYINPUT52,KEYINPUT53,G9,G75,G72,G69,G66,G63,G60,G6,G57,G54,G51,
G48,G45,G42,G39,G36,G33,G30,G3,G27,G24,G21,G18,G15,G12 );
input G953,
 G898, G224, G902, G952, G214, G900, G221, G110, G217, G119, G137, G128, G234, G472,
 G101, G210, G237, G125, G122, G113, G116, G469, G140, G227, G107, G104, G134, G131,
 G146, G475, G143, G478, KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9,
 KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
 KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37,
 KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51,
 KEYINPUT52, KEYINPUT53;
output G9, G75, G72, G69, G66, G63, G60, G6, G57, G54, G51, G48, G45, G42,
 G39, G36, G33, G30, G3, G27, G24, G21, G18, G15, G12;
XNOR_X1 U236 ( .A1(w1000), .A2(n211), .ZN(G9) );
NAND_X1 U237 ( .A1(n212), .A2(n213), .A3(n214), .ZN(G75) );
NOR_X1 U238 ( .A1(n215), .A2(G953), .A3(n216), .ZN(n214) );
NOR_X1 U239 ( .A1(n217), .A2(n218), .A3(n219), .A4(n220), .ZN(n216) );
NOR_X1 U240 ( .A1(n221), .A2(n222), .ZN(n217) );
NOR_X1 U241 ( .A1(n223), .A2(n224), .ZN(n222) );
NOR_X1 U242 ( .A1(n225), .A2(n226), .ZN(n223) );
NOR_X1 U243 ( .A1(n227), .A2(n228), .ZN(n221) );
NOR_X1 U244 ( .A1(n229), .A2(n230), .ZN(n227) );
NOR_X1 U245 ( .A1(n228), .A2(n231), .A3(n224), .ZN(n215) );
INV_X1 U246 ( .A1(n232), .ZN(n224) );
NOR_X1 U247 ( .A1(n233), .A2(n234), .ZN(n231) );
NOR_X1 U248 ( .A1(n218), .A2(n219), .ZN(n234) );
NOR_X1 U249 ( .A1(n235), .A2(n220), .ZN(n233) );
NOR_X1 U250 ( .A1(n236), .A2(n237), .ZN(n235) );
NOR_X1 U251 ( .A1(n238), .A2(n218), .ZN(n237) );
INV_X1 U252 ( .A1(n239), .ZN(n218) );
NOR_X1 U253 ( .A1(n240), .A2(n241), .ZN(n238) );
NOR_X1 U254 ( .A1(n242), .A2(n219), .ZN(n236) );
NOR_X1 U255 ( .A1(n243), .A2(n244), .ZN(n242) );
XOR_X1 U256 ( .A1(n245), .A2(n246), .ZN(w1004) );
XOR_X1 U257 ( .A1(n247), .A2(n248), .ZN(w1002) );
NOR_X1 U258 ( .A1(n249), .A2(n250), .ZN(w1005) );
NOR_X1 U259 ( .A1(n251), .A2(n252), .ZN(n249) );
NAND_X1 U260 ( .A1(n253), .A2(n254), .ZN(w1006) );
NAND_X1 U261 ( .A1(G953), .A2(n252), .ZN(n254) );
XOR_X1 U262 ( .A1(n255), .A2(n256), .ZN(n253) );
NAND_X1 U263 ( .A1(n250), .A2(n257), .ZN(w1003) );
XOR_X1 U264 ( .A1(n258), .A2(n259), .ZN(w1010) );
XOR_X1 U265 ( .A1(n260), .A2(n261), .ZN(w1008) );
NAND_X1 U266 ( .A1(n262), .A2(n263), .ZN(w1011) );
NAND_X1 U267 ( .A1(G953), .A2(n264), .ZN(n263) );
NAND_X1 U268 ( .A1(G953), .A2(n265), .ZN(n260) );
NAND_X1 U269 ( .A1(G898), .A2(G224), .ZN(n265) );
NOR_X1 U270 ( .A1(n212), .A2(G953), .ZN(w1009) );
NOR_X1 U271 ( .A1(n266), .A2(n267), .ZN(w1012) );
XNOR_X1 U272 ( .A1(n268), .A2(n269), .ZN(n267) );
NOR_X1 U273 ( .A1(n270), .A2(n271), .ZN(w1013) );
NOR_X1 U274 ( .A1(n266), .A2(n272), .ZN(w1014) );
XNOR_X1 U275 ( .A1(n273), .A2(n274), .ZN(n272) );
NOR_X1 U276 ( .A1(n275), .A2(n271), .ZN(w1015) );
NOR_X1 U277 ( .A1(n266), .A2(n276), .ZN(w1016) );
XNOR_X1 U278 ( .A1(n277), .A2(n278), .ZN(n276) );
NOR_X1 U279 ( .A1(n279), .A2(n271), .ZN(w1017) );
XNOR_X1 U280 ( .A1(w1018), .A2(n280), .ZN(G6) );
NOR_X1 U281 ( .A1(n266), .A2(n281), .ZN(w1020) );
XOR_X1 U282 ( .A1(n282), .A2(n283), .ZN(w1022) );
XOR_X1 U283 ( .A1(n284), .A2(n285), .ZN(w1021) );
NOR_X1 U284 ( .A1(n286), .A2(n271), .ZN(w1023) );
NOR_X1 U285 ( .A1(n266), .A2(n287), .ZN(w1024) );
XNOR_X1 U286 ( .A1(n288), .A2(n289), .ZN(n287) );
NOR_X1 U287 ( .A1(n290), .A2(n271), .ZN(w1025) );
NOR_X1 U288 ( .A1(n266), .A2(n291), .ZN(w1026) );
XNOR_X1 U289 ( .A1(n292), .A2(n293), .ZN(n291) );
NOR_X1 U290 ( .A1(n294), .A2(n271), .ZN(w1027) );
NAND_X1 U291 ( .A1(G902), .A2(n295), .ZN(n271) );
NAND_X1 U292 ( .A1(n212), .A2(n213), .ZN(n295) );
INV_X1 U293 ( .A1(n257), .ZN(n213) );
NAND_X1 U294 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(n257) );
NOR_X1 U295 ( .A1(n300), .A2(n301), .A3(n302), .A4(n303), .ZN(n299) );
NOR_X1 U296 ( .A1(n304), .A2(n305), .ZN(n298) );
AND_X1 U297 ( .A1(n306), .A2(n307), .ZN(n212) );
AND_X1 U298 ( .A1(n308), .A2(n309), .A3(n310), .A4(n311), .ZN(n307) );
AND_X1 U299 ( .A1(n312), .A2(n313), .A3(n211), .A4(n280), .ZN(n306) );
NAND_X1 U300 ( .A1(n239), .A2(n314), .A3(n230), .ZN(w1019) );
NAND_X1 U301 ( .A1(n239), .A2(n314), .A3(n229), .ZN(w1001) );
NOR_X1 U302 ( .A1(n250), .A2(G952), .ZN(n266) );
XNOR_X1 U303 ( .A1(w1028), .A2(n296), .ZN(G48) );
NAND_X1 U304 ( .A1(n230), .A2(n240), .A3(n315), .ZN(w1029) );
XNOR_X1 U305 ( .A1(w1030), .A2(n297), .ZN(G45) );
NAND_X1 U306 ( .A1(n316), .A2(n240), .A3(n317), .A4(n318), .ZN(w1031) );
XOR_X1 U307 ( .A1(w1032), .A2(n305), .ZN(G42) );
AND_X1 U308 ( .A1(n319), .A2(n225), .A3(n320), .ZN(w1033) );
XOR_X1 U309 ( .A1(w1034), .A2(n304), .ZN(G39) );
AND_X1 U310 ( .A1(n315), .A2(n232), .A3(n320), .ZN(w1035) );
XOR_X1 U311 ( .A1(w1036), .A2(n303), .ZN(G36) );
AND_X1 U312 ( .A1(n316), .A2(n229), .A3(n320), .ZN(w1037) );
XOR_X1 U313 ( .A1(w1038), .A2(n302), .ZN(G33) );
AND_X1 U314 ( .A1(n316), .A2(n230), .A3(n320), .ZN(w1039) );
INV_X1 U315 ( .A1(n219), .ZN(n320) );
NAND_X1 U316 ( .A1(n241), .A2(n321), .ZN(n219) );
NAND_X1 U317 ( .A1(G214), .A2(n322), .ZN(n321) );
AND_X1 U318 ( .A1(n225), .A2(n323), .A3(n243), .ZN(n316) );
XOR_X1 U319 ( .A1(w1040), .A2(n301), .ZN(G30) );
AND_X1 U320 ( .A1(n229), .A2(n240), .A3(n315), .ZN(w1041) );
AND_X1 U321 ( .A1(n225), .A2(n324), .A3(n325), .A4(n323), .ZN(n315) );
XNOR_X1 U322 ( .A1(w1042), .A2(n313), .ZN(G3) );
NAND_X1 U323 ( .A1(n232), .A2(n314), .A3(n243), .ZN(w1043) );
XOR_X1 U324 ( .A1(w1044), .A2(n300), .ZN(G27) );
AND_X1 U325 ( .A1(n326), .A2(n240), .A3(n319), .ZN(w1045) );
AND_X1 U326 ( .A1(n244), .A2(n230), .A3(n324), .A4(n323), .ZN(n319) );
NAND_X1 U327 ( .A1(n327), .A2(n220), .ZN(n323) );
NAND_X1 U328 ( .A1(n328), .A2(n252), .ZN(n327) );
INV_X1 U329 ( .A1(G900), .ZN(n252) );
XNOR_X1 U330 ( .A1(w1046), .A2(n312), .ZN(G24) );
NAND_X1 U331 ( .A1(n329), .A2(n239), .A3(n317), .A4(n318), .ZN(w1047) );
NOR_X1 U332 ( .A1(n325), .A2(n324), .ZN(n239) );
XNOR_X1 U333 ( .A1(w1048), .A2(n311), .ZN(G21) );
NAND_X1 U334 ( .A1(n329), .A2(n232), .A3(n324), .A4(n325), .ZN(w1049) );
XNOR_X1 U335 ( .A1(w1050), .A2(n310), .ZN(G18) );
NAND_X1 U336 ( .A1(n329), .A2(n229), .A3(n243), .ZN(w1051) );
NOR_X1 U337 ( .A1(n318), .A2(n330), .ZN(n229) );
XNOR_X1 U338 ( .A1(w1052), .A2(n309), .ZN(G15) );
NAND_X1 U339 ( .A1(n329), .A2(n230), .A3(n243), .ZN(w1053) );
NOR_X1 U340 ( .A1(n324), .A2(n244), .ZN(n243) );
AND_X1 U341 ( .A1(n330), .A2(n318), .ZN(n230) );
INV_X1 U342 ( .A1(n317), .ZN(n330) );
AND_X1 U343 ( .A1(n326), .A2(n331), .ZN(n329) );
INV_X1 U344 ( .A1(n228), .ZN(n326) );
NAND_X1 U345 ( .A1(n226), .A2(n332), .ZN(n228) );
NAND_X1 U346 ( .A1(G221), .A2(n333), .ZN(n332) );
XNOR_X1 U347 ( .A1(G110), .A2(n308), .ZN(G12) );
NAND_X1 U348 ( .A1(n232), .A2(n314), .A3(n244), .A4(n324), .ZN(n308) );
XOR_X1 U349 ( .A1(n334), .A2(n270), .ZN(n324) );
NAND_X1 U350 ( .A1(G217), .A2(n333), .ZN(n270) );
NAND_X1 U351 ( .A1(n268), .A2(n335), .ZN(n334) );
XNOR_X1 U352 ( .A1(n336), .A2(n337), .ZN(n268) );
XOR_X1 U353 ( .A1(G119), .A2(n338), .ZN(n337) );
XOR_X1 U354 ( .A1(G137), .A2(G128), .ZN(n338) );
XOR_X1 U355 ( .A1(n339), .A2(n340), .ZN(n336) );
XOR_X1 U356 ( .A1(G110), .A2(n341), .ZN(n340) );
AND_X1 U357 ( .A1(G221), .A2(n250), .A3(G234), .ZN(n341) );
INV_X1 U358 ( .A1(n325), .ZN(n244) );
XOR_X1 U359 ( .A1(n342), .A2(n286), .ZN(n325) );
INV_X1 U360 ( .A1(G472), .ZN(n286) );
NAND_X1 U361 ( .A1(n343), .A2(n335), .ZN(n342) );
XNOR_X1 U362 ( .A1(n284), .A2(n283), .ZN(n343) );
XNOR_X1 U363 ( .A1(n344), .A2(G101), .ZN(n283) );
NAND_X1 U364 ( .A1(G210), .A2(n345), .ZN(n344) );
XNOR_X1 U365 ( .A1(n255), .A2(n346), .ZN(n284) );
INV_X1 U366 ( .A1(n347), .ZN(n346) );
AND_X1 U367 ( .A1(n225), .A2(n331), .ZN(n314) );
AND_X1 U368 ( .A1(n240), .A2(n348), .ZN(n331) );
NAND_X1 U369 ( .A1(n349), .A2(n220), .ZN(n348) );
NAND_X1 U370 ( .A1(n350), .A2(n250), .A3(G952), .ZN(n220) );
NAND_X1 U371 ( .A1(n328), .A2(n264), .ZN(n349) );
INV_X1 U372 ( .A1(G898), .ZN(n264) );
AND_X1 U373 ( .A1(G902), .A2(n350), .A3(G953), .ZN(n328) );
NAND_X1 U374 ( .A1(G237), .A2(G234), .ZN(n350) );
NOR_X1 U375 ( .A1(n241), .A2(n351), .ZN(n240) );
AND_X1 U376 ( .A1(G214), .A2(n322), .ZN(n351) );
XNOR_X1 U377 ( .A1(n352), .A2(n294), .ZN(n241) );
NAND_X1 U378 ( .A1(G210), .A2(n322), .ZN(n294) );
NAND_X1 U379 ( .A1(n353), .A2(n335), .ZN(n322) );
INV_X1 U380 ( .A1(G237), .ZN(n353) );
NAND_X1 U381 ( .A1(n292), .A2(n335), .ZN(n352) );
XNOR_X1 U382 ( .A1(n354), .A2(n355), .ZN(n292) );
XOR_X1 U383 ( .A1(G125), .A2(n356), .ZN(n355) );
AND_X1 U384 ( .A1(n250), .A2(G224), .ZN(n356) );
XOR_X1 U385 ( .A1(n262), .A2(n357), .ZN(n354) );
XOR_X1 U386 ( .A1(n358), .A2(n359), .ZN(n262) );
XOR_X1 U387 ( .A1(G122), .A2(G110), .ZN(n359) );
XNOR_X1 U388 ( .A1(n347), .A2(n360), .ZN(n358) );
XOR_X1 U389 ( .A1(G113), .A2(n361), .ZN(n347) );
XOR_X1 U390 ( .A1(G119), .A2(G116), .ZN(n361) );
NOR_X1 U391 ( .A1(n226), .A2(n362), .ZN(n225) );
AND_X1 U392 ( .A1(G221), .A2(n333), .ZN(n362) );
NAND_X1 U393 ( .A1(G234), .A2(n335), .ZN(n333) );
XNOR_X1 U394 ( .A1(n363), .A2(n290), .ZN(n226) );
INV_X1 U395 ( .A1(G469), .ZN(n290) );
NAND_X1 U396 ( .A1(n288), .A2(n335), .ZN(n363) );
XNOR_X1 U397 ( .A1(n364), .A2(n365), .ZN(n288) );
XOR_X1 U398 ( .A1(n366), .A2(n367), .ZN(n365) );
XOR_X1 U399 ( .A1(G140), .A2(G110), .ZN(n367) );
NOR_X1 U400 ( .A1(G953), .A2(n251), .ZN(n366) );
INV_X1 U401 ( .A1(G227), .ZN(n251) );
XOR_X1 U402 ( .A1(n255), .A2(n360), .ZN(n364) );
XOR_X1 U403 ( .A1(G101), .A2(n368), .ZN(n360) );
XOR_X1 U404 ( .A1(G107), .A2(G104), .ZN(n368) );
XOR_X1 U405 ( .A1(n369), .A2(n370), .ZN(w1007) );
XOR_X1 U406 ( .A1(G137), .A2(G134), .ZN(n370) );
XNOR_X1 U407 ( .A1(n357), .A2(G131), .ZN(n369) );
XOR_X1 U408 ( .A1(G146), .A2(n371), .ZN(n357) );
NOR_X1 U409 ( .A1(n317), .A2(n318), .ZN(n232) );
XOR_X1 U410 ( .A1(n372), .A2(n279), .ZN(n318) );
INV_X1 U411 ( .A1(G475), .ZN(n279) );
NAND_X1 U412 ( .A1(n277), .A2(n335), .ZN(n372) );
XNOR_X1 U413 ( .A1(n373), .A2(n374), .ZN(n277) );
XOR_X1 U414 ( .A1(n375), .A2(n376), .ZN(n374) );
XOR_X1 U415 ( .A1(G122), .A2(G113), .ZN(n376) );
XNOR_X1 U416 ( .A1(n377), .A2(G131), .ZN(n375) );
INV_X1 U417 ( .A1(G143), .ZN(n377) );
XOR_X1 U418 ( .A1(n339), .A2(n378), .ZN(n373) );
XNOR_X1 U419 ( .A1(G104), .A2(n379), .ZN(n378) );
NAND_X1 U420 ( .A1(G214), .A2(n345), .ZN(n379) );
NOR_X1 U421 ( .A1(G953), .A2(G237), .ZN(n345) );
XNOR_X1 U422 ( .A1(G146), .A2(n256), .ZN(n339) );
XOR_X1 U423 ( .A1(G125), .A2(G140), .ZN(n256) );
XOR_X1 U424 ( .A1(n380), .A2(n275), .ZN(n317) );
INV_X1 U425 ( .A1(G478), .ZN(n275) );
NAND_X1 U426 ( .A1(n274), .A2(n335), .ZN(n380) );
INV_X1 U427 ( .A1(G902), .ZN(n335) );
NAND_X1 U428 ( .A1(n381), .A2(n382), .ZN(n274) );
NAND_X1 U429 ( .A1(n383), .A2(n384), .ZN(n382) );
NAND_X1 U430 ( .A1(G217), .A2(n250), .A3(G234), .ZN(n384) );
NAND_X1 U431 ( .A1(G217), .A2(n250), .A3(G234), .A4(n385), .ZN(n381) );
INV_X1 U432 ( .A1(n383), .ZN(n385) );
XNOR_X1 U433 ( .A1(n386), .A2(n387), .ZN(n383) );
XOR_X1 U434 ( .A1(G116), .A2(n388), .ZN(n387) );
XOR_X1 U435 ( .A1(G134), .A2(G122), .ZN(n388) );
XNOR_X1 U436 ( .A1(G107), .A2(n371), .ZN(n386) );
XOR_X1 U437 ( .A1(G128), .A2(G143), .ZN(n371) );
INV_X1 U438 ( .A1(G953), .ZN(n250) );
XOR_X1 X1000 ( .A1(G107), .A2(KEYINPUT0), .ZN(w1000) );
XNOR_X1 X1001 ( .A1(w1001), .A2(KEYINPUT1), .ZN(n211) );
XOR_X1 X1002 ( .A1(w1002), .A2(KEYINPUT2), .ZN(n246) );
XNOR_X1 X1003 ( .A1(w1003), .A2(KEYINPUT3), .ZN(n245) );
XOR_X1 X1004 ( .A1(w1004), .A2(KEYINPUT4), .ZN(G72) );
XNOR_X1 X1005 ( .A1(w1005), .A2(KEYINPUT5), .ZN(n248) );
XOR_X1 X1006 ( .A1(w1006), .A2(KEYINPUT6), .ZN(n247) );
XNOR_X1 X1007 ( .A1(w1007), .A2(KEYINPUT7), .ZN(n255) );
XOR_X1 X1008 ( .A1(w1008), .A2(KEYINPUT8), .ZN(n259) );
XNOR_X1 X1009 ( .A1(w1009), .A2(KEYINPUT9), .ZN(n258) );
XOR_X1 X1010 ( .A1(w1010), .A2(KEYINPUT10), .ZN(G69) );
XNOR_X1 X1011 ( .A1(w1011), .A2(KEYINPUT11), .ZN(n261) );
XOR_X1 X1012 ( .A1(w1012), .A2(KEYINPUT12), .ZN(G66) );
XNOR_X1 X1013 ( .A1(w1013), .A2(KEYINPUT13), .ZN(n269) );
XOR_X1 X1014 ( .A1(w1014), .A2(KEYINPUT14), .ZN(G63) );
XNOR_X1 X1015 ( .A1(w1015), .A2(KEYINPUT15), .ZN(n273) );
XOR_X1 X1016 ( .A1(w1016), .A2(KEYINPUT16), .ZN(G60) );
XNOR_X1 X1017 ( .A1(w1017), .A2(KEYINPUT17), .ZN(n278) );
XOR_X1 X1018 ( .A1(G104), .A2(KEYINPUT18), .ZN(w1018) );
XNOR_X1 X1019 ( .A1(w1019), .A2(KEYINPUT19), .ZN(n280) );
XOR_X1 X1020 ( .A1(w1020), .A2(KEYINPUT20), .ZN(G57) );
XNOR_X1 X1021 ( .A1(w1021), .A2(KEYINPUT21), .ZN(n282) );
XOR_X1 X1022 ( .A1(w1022), .A2(KEYINPUT22), .ZN(n281) );
XNOR_X1 X1023 ( .A1(w1023), .A2(KEYINPUT23), .ZN(n285) );
XOR_X1 X1024 ( .A1(w1024), .A2(KEYINPUT24), .ZN(G54) );
XNOR_X1 X1025 ( .A1(w1025), .A2(KEYINPUT25), .ZN(n289) );
XOR_X1 X1026 ( .A1(w1026), .A2(KEYINPUT26), .ZN(G51) );
XNOR_X1 X1027 ( .A1(w1027), .A2(KEYINPUT27), .ZN(n293) );
XOR_X1 X1028 ( .A1(G146), .A2(KEYINPUT28), .ZN(w1028) );
XNOR_X1 X1029 ( .A1(w1029), .A2(KEYINPUT29), .ZN(n296) );
XOR_X1 X1030 ( .A1(G143), .A2(KEYINPUT30), .ZN(w1030) );
XNOR_X1 X1031 ( .A1(w1031), .A2(KEYINPUT31), .ZN(n297) );
XOR_X1 X1032 ( .A1(G140), .A2(KEYINPUT32), .ZN(w1032) );
XNOR_X1 X1033 ( .A1(w1033), .A2(KEYINPUT33), .ZN(n305) );
XOR_X1 X1034 ( .A1(G137), .A2(KEYINPUT34), .ZN(w1034) );
XNOR_X1 X1035 ( .A1(w1035), .A2(KEYINPUT35), .ZN(n304) );
XOR_X1 X1036 ( .A1(G134), .A2(KEYINPUT36), .ZN(w1036) );
XNOR_X1 X1037 ( .A1(w1037), .A2(KEYINPUT37), .ZN(n303) );
XOR_X1 X1038 ( .A1(G131), .A2(KEYINPUT38), .ZN(w1038) );
XNOR_X1 X1039 ( .A1(w1039), .A2(KEYINPUT39), .ZN(n302) );
XOR_X1 X1040 ( .A1(G128), .A2(KEYINPUT40), .ZN(w1040) );
XNOR_X1 X1041 ( .A1(w1041), .A2(KEYINPUT41), .ZN(n301) );
XOR_X1 X1042 ( .A1(G101), .A2(KEYINPUT42), .ZN(w1042) );
XNOR_X1 X1043 ( .A1(w1043), .A2(KEYINPUT43), .ZN(n313) );
XOR_X1 X1044 ( .A1(G125), .A2(KEYINPUT44), .ZN(w1044) );
XNOR_X1 X1045 ( .A1(w1045), .A2(KEYINPUT45), .ZN(n300) );
XOR_X1 X1046 ( .A1(G122), .A2(KEYINPUT46), .ZN(w1046) );
XNOR_X1 X1047 ( .A1(w1047), .A2(KEYINPUT47), .ZN(n312) );
XOR_X1 X1048 ( .A1(G119), .A2(KEYINPUT48), .ZN(w1048) );
XNOR_X1 X1049 ( .A1(w1049), .A2(KEYINPUT49), .ZN(n311) );
XOR_X1 X1050 ( .A1(G116), .A2(KEYINPUT50), .ZN(w1050) );
XNOR_X1 X1051 ( .A1(w1051), .A2(KEYINPUT51), .ZN(n310) );
XOR_X1 X1052 ( .A1(G113), .A2(KEYINPUT52), .ZN(w1052) );
XNOR_X1 X1053 ( .A1(w1053), .A2(KEYINPUT53), .ZN(n309) );
